module carry_ripple_4bit(X, Y, C_in, S);
input [511:0] X;
input [511:0] Y;
input C_in;
output [512:0] S;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire _1889_;
wire _1890_;
wire _1891_;
wire _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire _1907_;
wire _1908_;
wire _1909_;
wire _1910_;
wire _1911_;
wire _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2053_;
wire _2054_;
wire _2055_;
wire _2056_;
wire _2057_;
wire _2058_;
wire _2059_;
wire _2060_;
wire _2061_;
wire _2062_;
wire _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
assign _1025_ = X[0] ^ Y[0];
assign _1026_ = X[0] & Y[0];
assign S[0] = _1025_ ^ C_in;
assign _1028_ = _1025_ & C_in;
assign _1029_ = _1026_ | _1028_;
assign _1030_ = X[1] ^ Y[1];
assign _1031_ = X[1] & Y[1];
assign S[1] = _1030_ ^ _1029_;
assign _1033_ = _1030_ & _1029_;
assign _1034_ = _1031_ | _1033_;
assign _1035_ = X[2] ^ Y[2];
assign _1036_ = X[2] & Y[2];
assign S[2] = _1035_ ^ _1034_;
assign _1038_ = _1035_ & _1034_;
assign _1039_ = _1036_ | _1038_;
assign _1040_ = X[3] ^ Y[3];
assign _1041_ = X[3] & Y[3];
assign S[3] = _1040_ ^ _1039_;
assign _1043_ = _1040_ & _1039_;
assign _1044_ = _1041_ | _1043_;
assign _1045_ = X[4] ^ Y[4];
assign _1046_ = X[4] & Y[4];
assign S[4] = _1045_ ^ _1044_;
assign _1048_ = _1045_ & _1044_;
assign _1049_ = _1046_ | _1048_;
assign _1050_ = X[5] ^ Y[5];
assign _1051_ = X[5] & Y[5];
assign S[5] = _1050_ ^ _1049_;
assign _1053_ = _1050_ & _1049_;
assign _1054_ = _1051_ | _1053_;
assign _1055_ = X[6] ^ Y[6];
assign _1056_ = X[6] & Y[6];
assign S[6] = _1055_ ^ _1054_;
assign _1058_ = _1055_ & _1054_;
assign _1059_ = _1056_ | _1058_;
assign _1060_ = X[7] ^ Y[7];
assign _1061_ = X[7] & Y[7];
assign S[7] = _1060_ ^ _1059_;
assign _1063_ = _1060_ & _1059_;
assign _1064_ = _1061_ | _1063_;
assign _1065_ = X[8] ^ Y[8];
assign _1066_ = X[8] & Y[8];
assign S[8] = _1065_ ^ _1064_;
assign _1068_ = _1065_ & _1064_;
assign _1069_ = _1066_ | _1068_;
assign _1070_ = X[9] ^ Y[9];
assign _1071_ = X[9] & Y[9];
assign S[9] = _1070_ ^ _1069_;
assign _1073_ = _1070_ & _1069_;
assign _1074_ = _1071_ | _1073_;
assign _1075_ = X[10] ^ Y[10];
assign _1076_ = X[10] & Y[10];
assign S[10] = _1075_ ^ _1074_;
assign _1078_ = _1075_ & _1074_;
assign _1079_ = _1076_ | _1078_;
assign _1080_ = X[11] ^ Y[11];
assign _1081_ = X[11] & Y[11];
assign S[11] = _1080_ ^ _1079_;
assign _1083_ = _1080_ & _1079_;
assign _1084_ = _1081_ | _1083_;
assign _1085_ = X[12] ^ Y[12];
assign _1086_ = X[12] & Y[12];
assign S[12] = _1085_ ^ _1084_;
assign _1088_ = _1085_ & _1084_;
assign _1089_ = _1086_ | _1088_;
assign _1090_ = X[13] ^ Y[13];
assign _1091_ = X[13] & Y[13];
assign S[13] = _1090_ ^ _1089_;
assign _1093_ = _1090_ & _1089_;
assign _1094_ = _1091_ | _1093_;
assign _1095_ = X[14] ^ Y[14];
assign _1096_ = X[14] & Y[14];
assign S[14] = _1095_ ^ _1094_;
assign _1098_ = _1095_ & _1094_;
assign _1099_ = _1096_ | _1098_;
assign _1100_ = X[15] ^ Y[15];
assign _1101_ = X[15] & Y[15];
assign S[15] = _1100_ ^ _1099_;
assign _1103_ = _1100_ & _1099_;
assign _1104_ = _1101_ | _1103_;
assign _1105_ = X[16] ^ Y[16];
assign _1106_ = X[16] & Y[16];
assign S[16] = _1105_ ^ _1104_;
assign _1108_ = _1105_ & _1104_;
assign _1109_ = _1106_ | _1108_;
assign _1110_ = X[17] ^ Y[17];
assign _1111_ = X[17] & Y[17];
assign S[17] = _1110_ ^ _1109_;
assign _1113_ = _1110_ & _1109_;
assign _1114_ = _1111_ | _1113_;
assign _1115_ = X[18] ^ Y[18];
assign _1116_ = X[18] & Y[18];
assign S[18] = _1115_ ^ _1114_;
assign _1118_ = _1115_ & _1114_;
assign _1119_ = _1116_ | _1118_;
assign _1120_ = X[19] ^ Y[19];
assign _1121_ = X[19] & Y[19];
assign S[19] = _1120_ ^ _1119_;
assign _1123_ = _1120_ & _1119_;
assign _1124_ = _1121_ | _1123_;
assign _1125_ = X[20] ^ Y[20];
assign _1126_ = X[20] & Y[20];
assign S[20] = _1125_ ^ _1124_;
assign _1128_ = _1125_ & _1124_;
assign _1129_ = _1126_ | _1128_;
assign _1130_ = X[21] ^ Y[21];
assign _1131_ = X[21] & Y[21];
assign S[21] = _1130_ ^ _1129_;
assign _1133_ = _1130_ & _1129_;
assign _1134_ = _1131_ | _1133_;
assign _1135_ = X[22] ^ Y[22];
assign _1136_ = X[22] & Y[22];
assign S[22] = _1135_ ^ _1134_;
assign _1138_ = _1135_ & _1134_;
assign _1139_ = _1136_ | _1138_;
assign _1140_ = X[23] ^ Y[23];
assign _1141_ = X[23] & Y[23];
assign S[23] = _1140_ ^ _1139_;
assign _1143_ = _1140_ & _1139_;
assign _1144_ = _1141_ | _1143_;
assign _1145_ = X[24] ^ Y[24];
assign _1146_ = X[24] & Y[24];
assign S[24] = _1145_ ^ _1144_;
assign _1148_ = _1145_ & _1144_;
assign _1149_ = _1146_ | _1148_;
assign _1150_ = X[25] ^ Y[25];
assign _1151_ = X[25] & Y[25];
assign S[25] = _1150_ ^ _1149_;
assign _1153_ = _1150_ & _1149_;
assign _1154_ = _1151_ | _1153_;
assign _1155_ = X[26] ^ Y[26];
assign _1156_ = X[26] & Y[26];
assign S[26] = _1155_ ^ _1154_;
assign _1158_ = _1155_ & _1154_;
assign _1159_ = _1156_ | _1158_;
assign _1160_ = X[27] ^ Y[27];
assign _1161_ = X[27] & Y[27];
assign S[27] = _1160_ ^ _1159_;
assign _1163_ = _1160_ & _1159_;
assign _1164_ = _1161_ | _1163_;
assign _1165_ = X[28] ^ Y[28];
assign _1166_ = X[28] & Y[28];
assign S[28] = _1165_ ^ _1164_;
assign _1168_ = _1165_ & _1164_;
assign _1169_ = _1166_ | _1168_;
assign _1170_ = X[29] ^ Y[29];
assign _1171_ = X[29] & Y[29];
assign S[29] = _1170_ ^ _1169_;
assign _1173_ = _1170_ & _1169_;
assign _1174_ = _1171_ | _1173_;
assign _1175_ = X[30] ^ Y[30];
assign _1176_ = X[30] & Y[30];
assign S[30] = _1175_ ^ _1174_;
assign _1178_ = _1175_ & _1174_;
assign _1179_ = _1176_ | _1178_;
assign _1180_ = X[31] ^ Y[31];
assign _1181_ = X[31] & Y[31];
assign S[31] = _1180_ ^ _1179_;
assign _1183_ = _1180_ & _1179_;
assign _1184_ = _1181_ | _1183_;
assign _1185_ = X[32] ^ Y[32];
assign _1186_ = X[32] & Y[32];
assign S[32] = _1185_ ^ _1184_;
assign _1188_ = _1185_ & _1184_;
assign _1189_ = _1186_ | _1188_;
assign _1190_ = X[33] ^ Y[33];
assign _1191_ = X[33] & Y[33];
assign S[33] = _1190_ ^ _1189_;
assign _1193_ = _1190_ & _1189_;
assign _1194_ = _1191_ | _1193_;
assign _1195_ = X[34] ^ Y[34];
assign _1196_ = X[34] & Y[34];
assign S[34] = _1195_ ^ _1194_;
assign _1198_ = _1195_ & _1194_;
assign _1199_ = _1196_ | _1198_;
assign _1200_ = X[35] ^ Y[35];
assign _1201_ = X[35] & Y[35];
assign S[35] = _1200_ ^ _1199_;
assign _1203_ = _1200_ & _1199_;
assign _1204_ = _1201_ | _1203_;
assign _1205_ = X[36] ^ Y[36];
assign _1206_ = X[36] & Y[36];
assign S[36] = _1205_ ^ _1204_;
assign _1208_ = _1205_ & _1204_;
assign _1209_ = _1206_ | _1208_;
assign _1210_ = X[37] ^ Y[37];
assign _1211_ = X[37] & Y[37];
assign S[37] = _1210_ ^ _1209_;
assign _1213_ = _1210_ & _1209_;
assign _1214_ = _1211_ | _1213_;
assign _1215_ = X[38] ^ Y[38];
assign _1216_ = X[38] & Y[38];
assign S[38] = _1215_ ^ _1214_;
assign _1218_ = _1215_ & _1214_;
assign _1219_ = _1216_ | _1218_;
assign _1220_ = X[39] ^ Y[39];
assign _1221_ = X[39] & Y[39];
assign S[39] = _1220_ ^ _1219_;
assign _1223_ = _1220_ & _1219_;
assign _1224_ = _1221_ | _1223_;
assign _1225_ = X[40] ^ Y[40];
assign _1226_ = X[40] & Y[40];
assign S[40] = _1225_ ^ _1224_;
assign _1228_ = _1225_ & _1224_;
assign _1229_ = _1226_ | _1228_;
assign _1230_ = X[41] ^ Y[41];
assign _1231_ = X[41] & Y[41];
assign S[41] = _1230_ ^ _1229_;
assign _1233_ = _1230_ & _1229_;
assign _1234_ = _1231_ | _1233_;
assign _1235_ = X[42] ^ Y[42];
assign _1236_ = X[42] & Y[42];
assign S[42] = _1235_ ^ _1234_;
assign _1238_ = _1235_ & _1234_;
assign _1239_ = _1236_ | _1238_;
assign _1240_ = X[43] ^ Y[43];
assign _1241_ = X[43] & Y[43];
assign S[43] = _1240_ ^ _1239_;
assign _1243_ = _1240_ & _1239_;
assign _1244_ = _1241_ | _1243_;
assign _1245_ = X[44] ^ Y[44];
assign _1246_ = X[44] & Y[44];
assign S[44] = _1245_ ^ _1244_;
assign _1248_ = _1245_ & _1244_;
assign _1249_ = _1246_ | _1248_;
assign _1250_ = X[45] ^ Y[45];
assign _1251_ = X[45] & Y[45];
assign S[45] = _1250_ ^ _1249_;
assign _1253_ = _1250_ & _1249_;
assign _1254_ = _1251_ | _1253_;
assign _1255_ = X[46] ^ Y[46];
assign _1256_ = X[46] & Y[46];
assign S[46] = _1255_ ^ _1254_;
assign _1258_ = _1255_ & _1254_;
assign _1259_ = _1256_ | _1258_;
assign _1260_ = X[47] ^ Y[47];
assign _1261_ = X[47] & Y[47];
assign S[47] = _1260_ ^ _1259_;
assign _1263_ = _1260_ & _1259_;
assign _1264_ = _1261_ | _1263_;
assign _1265_ = X[48] ^ Y[48];
assign _1266_ = X[48] & Y[48];
assign S[48] = _1265_ ^ _1264_;
assign _1268_ = _1265_ & _1264_;
assign _1269_ = _1266_ | _1268_;
assign _1270_ = X[49] ^ Y[49];
assign _1271_ = X[49] & Y[49];
assign S[49] = _1270_ ^ _1269_;
assign _1273_ = _1270_ & _1269_;
assign _1274_ = _1271_ | _1273_;
assign _1275_ = X[50] ^ Y[50];
assign _1276_ = X[50] & Y[50];
assign S[50] = _1275_ ^ _1274_;
assign _1278_ = _1275_ & _1274_;
assign _1279_ = _1276_ | _1278_;
assign _1280_ = X[51] ^ Y[51];
assign _1281_ = X[51] & Y[51];
assign S[51] = _1280_ ^ _1279_;
assign _1283_ = _1280_ & _1279_;
assign _1284_ = _1281_ | _1283_;
assign _1285_ = X[52] ^ Y[52];
assign _1286_ = X[52] & Y[52];
assign S[52] = _1285_ ^ _1284_;
assign _1288_ = _1285_ & _1284_;
assign _1289_ = _1286_ | _1288_;
assign _1290_ = X[53] ^ Y[53];
assign _1291_ = X[53] & Y[53];
assign S[53] = _1290_ ^ _1289_;
assign _1293_ = _1290_ & _1289_;
assign _1294_ = _1291_ | _1293_;
assign _1295_ = X[54] ^ Y[54];
assign _1296_ = X[54] & Y[54];
assign S[54] = _1295_ ^ _1294_;
assign _1298_ = _1295_ & _1294_;
assign _1299_ = _1296_ | _1298_;
assign _1300_ = X[55] ^ Y[55];
assign _1301_ = X[55] & Y[55];
assign S[55] = _1300_ ^ _1299_;
assign _1303_ = _1300_ & _1299_;
assign _1304_ = _1301_ | _1303_;
assign _1305_ = X[56] ^ Y[56];
assign _1306_ = X[56] & Y[56];
assign S[56] = _1305_ ^ _1304_;
assign _1308_ = _1305_ & _1304_;
assign _1309_ = _1306_ | _1308_;
assign _1310_ = X[57] ^ Y[57];
assign _1311_ = X[57] & Y[57];
assign S[57] = _1310_ ^ _1309_;
assign _1313_ = _1310_ & _1309_;
assign _1314_ = _1311_ | _1313_;
assign _1315_ = X[58] ^ Y[58];
assign _1316_ = X[58] & Y[58];
assign S[58] = _1315_ ^ _1314_;
assign _1318_ = _1315_ & _1314_;
assign _1319_ = _1316_ | _1318_;
assign _1320_ = X[59] ^ Y[59];
assign _1321_ = X[59] & Y[59];
assign S[59] = _1320_ ^ _1319_;
assign _1323_ = _1320_ & _1319_;
assign _1324_ = _1321_ | _1323_;
assign _1325_ = X[60] ^ Y[60];
assign _1326_ = X[60] & Y[60];
assign S[60] = _1325_ ^ _1324_;
assign _1328_ = _1325_ & _1324_;
assign _1329_ = _1326_ | _1328_;
assign _1330_ = X[61] ^ Y[61];
assign _1331_ = X[61] & Y[61];
assign S[61] = _1330_ ^ _1329_;
assign _1333_ = _1330_ & _1329_;
assign _1334_ = _1331_ | _1333_;
assign _1335_ = X[62] ^ Y[62];
assign _1336_ = X[62] & Y[62];
assign S[62] = _1335_ ^ _1334_;
assign _1338_ = _1335_ & _1334_;
assign _1339_ = _1336_ | _1338_;
assign _1340_ = X[63] ^ Y[63];
assign _1341_ = X[63] & Y[63];
assign S[63] = _1340_ ^ _1339_;
assign _1343_ = _1340_ & _1339_;
assign _1344_ = _1341_ | _1343_;
assign _1345_ = X[64] ^ Y[64];
assign _1346_ = X[64] & Y[64];
assign S[64] = _1345_ ^ _1344_;
assign _1348_ = _1345_ & _1344_;
assign _1349_ = _1346_ | _1348_;
assign _1350_ = X[65] ^ Y[65];
assign _1351_ = X[65] & Y[65];
assign S[65] = _1350_ ^ _1349_;
assign _1353_ = _1350_ & _1349_;
assign _1354_ = _1351_ | _1353_;
assign _1355_ = X[66] ^ Y[66];
assign _1356_ = X[66] & Y[66];
assign S[66] = _1355_ ^ _1354_;
assign _1358_ = _1355_ & _1354_;
assign _1359_ = _1356_ | _1358_;
assign _1360_ = X[67] ^ Y[67];
assign _1361_ = X[67] & Y[67];
assign S[67] = _1360_ ^ _1359_;
assign _1363_ = _1360_ & _1359_;
assign _1364_ = _1361_ | _1363_;
assign _1365_ = X[68] ^ Y[68];
assign _1366_ = X[68] & Y[68];
assign S[68] = _1365_ ^ _1364_;
assign _1368_ = _1365_ & _1364_;
assign _1369_ = _1366_ | _1368_;
assign _1370_ = X[69] ^ Y[69];
assign _1371_ = X[69] & Y[69];
assign S[69] = _1370_ ^ _1369_;
assign _1373_ = _1370_ & _1369_;
assign _1374_ = _1371_ | _1373_;
assign _1375_ = X[70] ^ Y[70];
assign _1376_ = X[70] & Y[70];
assign S[70] = _1375_ ^ _1374_;
assign _1378_ = _1375_ & _1374_;
assign _1379_ = _1376_ | _1378_;
assign _1380_ = X[71] ^ Y[71];
assign _1381_ = X[71] & Y[71];
assign S[71] = _1380_ ^ _1379_;
assign _1383_ = _1380_ & _1379_;
assign _1384_ = _1381_ | _1383_;
assign _1385_ = X[72] ^ Y[72];
assign _1386_ = X[72] & Y[72];
assign S[72] = _1385_ ^ _1384_;
assign _1388_ = _1385_ & _1384_;
assign _1389_ = _1386_ | _1388_;
assign _1390_ = X[73] ^ Y[73];
assign _1391_ = X[73] & Y[73];
assign S[73] = _1390_ ^ _1389_;
assign _1393_ = _1390_ & _1389_;
assign _1394_ = _1391_ | _1393_;
assign _1395_ = X[74] ^ Y[74];
assign _1396_ = X[74] & Y[74];
assign S[74] = _1395_ ^ _1394_;
assign _1398_ = _1395_ & _1394_;
assign _1399_ = _1396_ | _1398_;
assign _1400_ = X[75] ^ Y[75];
assign _1401_ = X[75] & Y[75];
assign S[75] = _1400_ ^ _1399_;
assign _1403_ = _1400_ & _1399_;
assign _1404_ = _1401_ | _1403_;
assign _1405_ = X[76] ^ Y[76];
assign _1406_ = X[76] & Y[76];
assign S[76] = _1405_ ^ _1404_;
assign _1408_ = _1405_ & _1404_;
assign _1409_ = _1406_ | _1408_;
assign _1410_ = X[77] ^ Y[77];
assign _1411_ = X[77] & Y[77];
assign S[77] = _1410_ ^ _1409_;
assign _1413_ = _1410_ & _1409_;
assign _1414_ = _1411_ | _1413_;
assign _1415_ = X[78] ^ Y[78];
assign _1416_ = X[78] & Y[78];
assign S[78] = _1415_ ^ _1414_;
assign _1418_ = _1415_ & _1414_;
assign _1419_ = _1416_ | _1418_;
assign _1420_ = X[79] ^ Y[79];
assign _1421_ = X[79] & Y[79];
assign S[79] = _1420_ ^ _1419_;
assign _1423_ = _1420_ & _1419_;
assign _1424_ = _1421_ | _1423_;
assign _1425_ = X[80] ^ Y[80];
assign _1426_ = X[80] & Y[80];
assign S[80] = _1425_ ^ _1424_;
assign _1428_ = _1425_ & _1424_;
assign _1429_ = _1426_ | _1428_;
assign _1430_ = X[81] ^ Y[81];
assign _1431_ = X[81] & Y[81];
assign S[81] = _1430_ ^ _1429_;
assign _1433_ = _1430_ & _1429_;
assign _1434_ = _1431_ | _1433_;
assign _1435_ = X[82] ^ Y[82];
assign _1436_ = X[82] & Y[82];
assign S[82] = _1435_ ^ _1434_;
assign _1438_ = _1435_ & _1434_;
assign _1439_ = _1436_ | _1438_;
assign _1440_ = X[83] ^ Y[83];
assign _1441_ = X[83] & Y[83];
assign S[83] = _1440_ ^ _1439_;
assign _1443_ = _1440_ & _1439_;
assign _1444_ = _1441_ | _1443_;
assign _1445_ = X[84] ^ Y[84];
assign _1446_ = X[84] & Y[84];
assign S[84] = _1445_ ^ _1444_;
assign _1448_ = _1445_ & _1444_;
assign _1449_ = _1446_ | _1448_;
assign _1450_ = X[85] ^ Y[85];
assign _1451_ = X[85] & Y[85];
assign S[85] = _1450_ ^ _1449_;
assign _1453_ = _1450_ & _1449_;
assign _1454_ = _1451_ | _1453_;
assign _1455_ = X[86] ^ Y[86];
assign _1456_ = X[86] & Y[86];
assign S[86] = _1455_ ^ _1454_;
assign _1458_ = _1455_ & _1454_;
assign _1459_ = _1456_ | _1458_;
assign _1460_ = X[87] ^ Y[87];
assign _1461_ = X[87] & Y[87];
assign S[87] = _1460_ ^ _1459_;
assign _1463_ = _1460_ & _1459_;
assign _1464_ = _1461_ | _1463_;
assign _1465_ = X[88] ^ Y[88];
assign _1466_ = X[88] & Y[88];
assign S[88] = _1465_ ^ _1464_;
assign _1468_ = _1465_ & _1464_;
assign _1469_ = _1466_ | _1468_;
assign _1470_ = X[89] ^ Y[89];
assign _1471_ = X[89] & Y[89];
assign S[89] = _1470_ ^ _1469_;
assign _1473_ = _1470_ & _1469_;
assign _1474_ = _1471_ | _1473_;
assign _1475_ = X[90] ^ Y[90];
assign _1476_ = X[90] & Y[90];
assign S[90] = _1475_ ^ _1474_;
assign _1478_ = _1475_ & _1474_;
assign _1479_ = _1476_ | _1478_;
assign _1480_ = X[91] ^ Y[91];
assign _1481_ = X[91] & Y[91];
assign S[91] = _1480_ ^ _1479_;
assign _1483_ = _1480_ & _1479_;
assign _1484_ = _1481_ | _1483_;
assign _1485_ = X[92] ^ Y[92];
assign _1486_ = X[92] & Y[92];
assign S[92] = _1485_ ^ _1484_;
assign _1488_ = _1485_ & _1484_;
assign _1489_ = _1486_ | _1488_;
assign _1490_ = X[93] ^ Y[93];
assign _1491_ = X[93] & Y[93];
assign S[93] = _1490_ ^ _1489_;
assign _1493_ = _1490_ & _1489_;
assign _1494_ = _1491_ | _1493_;
assign _1495_ = X[94] ^ Y[94];
assign _1496_ = X[94] & Y[94];
assign S[94] = _1495_ ^ _1494_;
assign _1498_ = _1495_ & _1494_;
assign _1499_ = _1496_ | _1498_;
assign _1500_ = X[95] ^ Y[95];
assign _1501_ = X[95] & Y[95];
assign S[95] = _1500_ ^ _1499_;
assign _1503_ = _1500_ & _1499_;
assign _1504_ = _1501_ | _1503_;
assign _1505_ = X[96] ^ Y[96];
assign _1506_ = X[96] & Y[96];
assign S[96] = _1505_ ^ _1504_;
assign _1508_ = _1505_ & _1504_;
assign _1509_ = _1506_ | _1508_;
assign _1510_ = X[97] ^ Y[97];
assign _1511_ = X[97] & Y[97];
assign S[97] = _1510_ ^ _1509_;
assign _1513_ = _1510_ & _1509_;
assign _1514_ = _1511_ | _1513_;
assign _1515_ = X[98] ^ Y[98];
assign _1516_ = X[98] & Y[98];
assign S[98] = _1515_ ^ _1514_;
assign _1518_ = _1515_ & _1514_;
assign _1519_ = _1516_ | _1518_;
assign _1520_ = X[99] ^ Y[99];
assign _1521_ = X[99] & Y[99];
assign S[99] = _1520_ ^ _1519_;
assign _1523_ = _1520_ & _1519_;
assign _1524_ = _1521_ | _1523_;
assign _1525_ = X[100] ^ Y[100];
assign _1526_ = X[100] & Y[100];
assign S[100] = _1525_ ^ _1524_;
assign _1528_ = _1525_ & _1524_;
assign _1529_ = _1526_ | _1528_;
assign _1530_ = X[101] ^ Y[101];
assign _1531_ = X[101] & Y[101];
assign S[101] = _1530_ ^ _1529_;
assign _1533_ = _1530_ & _1529_;
assign _1534_ = _1531_ | _1533_;
assign _1535_ = X[102] ^ Y[102];
assign _1536_ = X[102] & Y[102];
assign S[102] = _1535_ ^ _1534_;
assign _1538_ = _1535_ & _1534_;
assign _1539_ = _1536_ | _1538_;
assign _1540_ = X[103] ^ Y[103];
assign _1541_ = X[103] & Y[103];
assign S[103] = _1540_ ^ _1539_;
assign _1543_ = _1540_ & _1539_;
assign _1544_ = _1541_ | _1543_;
assign _1545_ = X[104] ^ Y[104];
assign _1546_ = X[104] & Y[104];
assign S[104] = _1545_ ^ _1544_;
assign _1548_ = _1545_ & _1544_;
assign _1549_ = _1546_ | _1548_;
assign _1550_ = X[105] ^ Y[105];
assign _1551_ = X[105] & Y[105];
assign S[105] = _1550_ ^ _1549_;
assign _1553_ = _1550_ & _1549_;
assign _1554_ = _1551_ | _1553_;
assign _1555_ = X[106] ^ Y[106];
assign _1556_ = X[106] & Y[106];
assign S[106] = _1555_ ^ _1554_;
assign _1558_ = _1555_ & _1554_;
assign _1559_ = _1556_ | _1558_;
assign _1560_ = X[107] ^ Y[107];
assign _1561_ = X[107] & Y[107];
assign S[107] = _1560_ ^ _1559_;
assign _1563_ = _1560_ & _1559_;
assign _1564_ = _1561_ | _1563_;
assign _1565_ = X[108] ^ Y[108];
assign _1566_ = X[108] & Y[108];
assign S[108] = _1565_ ^ _1564_;
assign _1568_ = _1565_ & _1564_;
assign _1569_ = _1566_ | _1568_;
assign _1570_ = X[109] ^ Y[109];
assign _1571_ = X[109] & Y[109];
assign S[109] = _1570_ ^ _1569_;
assign _1573_ = _1570_ & _1569_;
assign _1574_ = _1571_ | _1573_;
assign _1575_ = X[110] ^ Y[110];
assign _1576_ = X[110] & Y[110];
assign S[110] = _1575_ ^ _1574_;
assign _1578_ = _1575_ & _1574_;
assign _1579_ = _1576_ | _1578_;
assign _1580_ = X[111] ^ Y[111];
assign _1581_ = X[111] & Y[111];
assign S[111] = _1580_ ^ _1579_;
assign _1583_ = _1580_ & _1579_;
assign _1584_ = _1581_ | _1583_;
assign _1585_ = X[112] ^ Y[112];
assign _1586_ = X[112] & Y[112];
assign S[112] = _1585_ ^ _1584_;
assign _1588_ = _1585_ & _1584_;
assign _1589_ = _1586_ | _1588_;
assign _1590_ = X[113] ^ Y[113];
assign _1591_ = X[113] & Y[113];
assign S[113] = _1590_ ^ _1589_;
assign _1593_ = _1590_ & _1589_;
assign _1594_ = _1591_ | _1593_;
assign _1595_ = X[114] ^ Y[114];
assign _1596_ = X[114] & Y[114];
assign S[114] = _1595_ ^ _1594_;
assign _1598_ = _1595_ & _1594_;
assign _1599_ = _1596_ | _1598_;
assign _1600_ = X[115] ^ Y[115];
assign _1601_ = X[115] & Y[115];
assign S[115] = _1600_ ^ _1599_;
assign _1603_ = _1600_ & _1599_;
assign _1604_ = _1601_ | _1603_;
assign _1605_ = X[116] ^ Y[116];
assign _1606_ = X[116] & Y[116];
assign S[116] = _1605_ ^ _1604_;
assign _1608_ = _1605_ & _1604_;
assign _1609_ = _1606_ | _1608_;
assign _1610_ = X[117] ^ Y[117];
assign _1611_ = X[117] & Y[117];
assign S[117] = _1610_ ^ _1609_;
assign _1613_ = _1610_ & _1609_;
assign _1614_ = _1611_ | _1613_;
assign _1615_ = X[118] ^ Y[118];
assign _1616_ = X[118] & Y[118];
assign S[118] = _1615_ ^ _1614_;
assign _1618_ = _1615_ & _1614_;
assign _1619_ = _1616_ | _1618_;
assign _1620_ = X[119] ^ Y[119];
assign _1621_ = X[119] & Y[119];
assign S[119] = _1620_ ^ _1619_;
assign _1623_ = _1620_ & _1619_;
assign _1624_ = _1621_ | _1623_;
assign _1625_ = X[120] ^ Y[120];
assign _1626_ = X[120] & Y[120];
assign S[120] = _1625_ ^ _1624_;
assign _1628_ = _1625_ & _1624_;
assign _1629_ = _1626_ | _1628_;
assign _1630_ = X[121] ^ Y[121];
assign _1631_ = X[121] & Y[121];
assign S[121] = _1630_ ^ _1629_;
assign _1633_ = _1630_ & _1629_;
assign _1634_ = _1631_ | _1633_;
assign _1635_ = X[122] ^ Y[122];
assign _1636_ = X[122] & Y[122];
assign S[122] = _1635_ ^ _1634_;
assign _1638_ = _1635_ & _1634_;
assign _1639_ = _1636_ | _1638_;
assign _1640_ = X[123] ^ Y[123];
assign _1641_ = X[123] & Y[123];
assign S[123] = _1640_ ^ _1639_;
assign _1643_ = _1640_ & _1639_;
assign _1644_ = _1641_ | _1643_;
assign _1645_ = X[124] ^ Y[124];
assign _1646_ = X[124] & Y[124];
assign S[124] = _1645_ ^ _1644_;
assign _1648_ = _1645_ & _1644_;
assign _1649_ = _1646_ | _1648_;
assign _1650_ = X[125] ^ Y[125];
assign _1651_ = X[125] & Y[125];
assign S[125] = _1650_ ^ _1649_;
assign _1653_ = _1650_ & _1649_;
assign _1654_ = _1651_ | _1653_;
assign _1655_ = X[126] ^ Y[126];
assign _1656_ = X[126] & Y[126];
assign S[126] = _1655_ ^ _1654_;
assign _1658_ = _1655_ & _1654_;
assign _1659_ = _1656_ | _1658_;
assign _1660_ = X[127] ^ Y[127];
assign _1661_ = X[127] & Y[127];
assign S[127] = _1660_ ^ _1659_;
assign _1663_ = _1660_ & _1659_;
assign _1664_ = _1661_ | _1663_;
assign _1665_ = X[128] ^ Y[128];
assign _1666_ = X[128] & Y[128];
assign S[128] = _1665_ ^ _1664_;
assign _1668_ = _1665_ & _1664_;
assign _1669_ = _1666_ | _1668_;
assign _1670_ = X[129] ^ Y[129];
assign _1671_ = X[129] & Y[129];
assign S[129] = _1670_ ^ _1669_;
assign _1673_ = _1670_ & _1669_;
assign _1674_ = _1671_ | _1673_;
assign _1675_ = X[130] ^ Y[130];
assign _1676_ = X[130] & Y[130];
assign S[130] = _1675_ ^ _1674_;
assign _1678_ = _1675_ & _1674_;
assign _1679_ = _1676_ | _1678_;
assign _1680_ = X[131] ^ Y[131];
assign _1681_ = X[131] & Y[131];
assign S[131] = _1680_ ^ _1679_;
assign _1683_ = _1680_ & _1679_;
assign _1684_ = _1681_ | _1683_;
assign _1685_ = X[132] ^ Y[132];
assign _1686_ = X[132] & Y[132];
assign S[132] = _1685_ ^ _1684_;
assign _1688_ = _1685_ & _1684_;
assign _1689_ = _1686_ | _1688_;
assign _1690_ = X[133] ^ Y[133];
assign _1691_ = X[133] & Y[133];
assign S[133] = _1690_ ^ _1689_;
assign _1693_ = _1690_ & _1689_;
assign _1694_ = _1691_ | _1693_;
assign _1695_ = X[134] ^ Y[134];
assign _1696_ = X[134] & Y[134];
assign S[134] = _1695_ ^ _1694_;
assign _1698_ = _1695_ & _1694_;
assign _1699_ = _1696_ | _1698_;
assign _1700_ = X[135] ^ Y[135];
assign _1701_ = X[135] & Y[135];
assign S[135] = _1700_ ^ _1699_;
assign _1703_ = _1700_ & _1699_;
assign _1704_ = _1701_ | _1703_;
assign _1705_ = X[136] ^ Y[136];
assign _1706_ = X[136] & Y[136];
assign S[136] = _1705_ ^ _1704_;
assign _1708_ = _1705_ & _1704_;
assign _1709_ = _1706_ | _1708_;
assign _1710_ = X[137] ^ Y[137];
assign _1711_ = X[137] & Y[137];
assign S[137] = _1710_ ^ _1709_;
assign _1713_ = _1710_ & _1709_;
assign _1714_ = _1711_ | _1713_;
assign _1715_ = X[138] ^ Y[138];
assign _1716_ = X[138] & Y[138];
assign S[138] = _1715_ ^ _1714_;
assign _1718_ = _1715_ & _1714_;
assign _1719_ = _1716_ | _1718_;
assign _1720_ = X[139] ^ Y[139];
assign _1721_ = X[139] & Y[139];
assign S[139] = _1720_ ^ _1719_;
assign _1723_ = _1720_ & _1719_;
assign _1724_ = _1721_ | _1723_;
assign _1725_ = X[140] ^ Y[140];
assign _1726_ = X[140] & Y[140];
assign S[140] = _1725_ ^ _1724_;
assign _1728_ = _1725_ & _1724_;
assign _1729_ = _1726_ | _1728_;
assign _1730_ = X[141] ^ Y[141];
assign _1731_ = X[141] & Y[141];
assign S[141] = _1730_ ^ _1729_;
assign _1733_ = _1730_ & _1729_;
assign _1734_ = _1731_ | _1733_;
assign _1735_ = X[142] ^ Y[142];
assign _1736_ = X[142] & Y[142];
assign S[142] = _1735_ ^ _1734_;
assign _1738_ = _1735_ & _1734_;
assign _1739_ = _1736_ | _1738_;
assign _1740_ = X[143] ^ Y[143];
assign _1741_ = X[143] & Y[143];
assign S[143] = _1740_ ^ _1739_;
assign _1743_ = _1740_ & _1739_;
assign _1744_ = _1741_ | _1743_;
assign _1745_ = X[144] ^ Y[144];
assign _1746_ = X[144] & Y[144];
assign S[144] = _1745_ ^ _1744_;
assign _1748_ = _1745_ & _1744_;
assign _1749_ = _1746_ | _1748_;
assign _1750_ = X[145] ^ Y[145];
assign _1751_ = X[145] & Y[145];
assign S[145] = _1750_ ^ _1749_;
assign _1753_ = _1750_ & _1749_;
assign _1754_ = _1751_ | _1753_;
assign _1755_ = X[146] ^ Y[146];
assign _1756_ = X[146] & Y[146];
assign S[146] = _1755_ ^ _1754_;
assign _1758_ = _1755_ & _1754_;
assign _1759_ = _1756_ | _1758_;
assign _1760_ = X[147] ^ Y[147];
assign _1761_ = X[147] & Y[147];
assign S[147] = _1760_ ^ _1759_;
assign _1763_ = _1760_ & _1759_;
assign _1764_ = _1761_ | _1763_;
assign _1765_ = X[148] ^ Y[148];
assign _1766_ = X[148] & Y[148];
assign S[148] = _1765_ ^ _1764_;
assign _1768_ = _1765_ & _1764_;
assign _1769_ = _1766_ | _1768_;
assign _1770_ = X[149] ^ Y[149];
assign _1771_ = X[149] & Y[149];
assign S[149] = _1770_ ^ _1769_;
assign _1773_ = _1770_ & _1769_;
assign _1774_ = _1771_ | _1773_;
assign _1775_ = X[150] ^ Y[150];
assign _1776_ = X[150] & Y[150];
assign S[150] = _1775_ ^ _1774_;
assign _1778_ = _1775_ & _1774_;
assign _1779_ = _1776_ | _1778_;
assign _1780_ = X[151] ^ Y[151];
assign _1781_ = X[151] & Y[151];
assign S[151] = _1780_ ^ _1779_;
assign _1783_ = _1780_ & _1779_;
assign _1784_ = _1781_ | _1783_;
assign _1785_ = X[152] ^ Y[152];
assign _1786_ = X[152] & Y[152];
assign S[152] = _1785_ ^ _1784_;
assign _1788_ = _1785_ & _1784_;
assign _1789_ = _1786_ | _1788_;
assign _1790_ = X[153] ^ Y[153];
assign _1791_ = X[153] & Y[153];
assign S[153] = _1790_ ^ _1789_;
assign _1793_ = _1790_ & _1789_;
assign _1794_ = _1791_ | _1793_;
assign _1795_ = X[154] ^ Y[154];
assign _1796_ = X[154] & Y[154];
assign S[154] = _1795_ ^ _1794_;
assign _1798_ = _1795_ & _1794_;
assign _1799_ = _1796_ | _1798_;
assign _1800_ = X[155] ^ Y[155];
assign _1801_ = X[155] & Y[155];
assign S[155] = _1800_ ^ _1799_;
assign _1803_ = _1800_ & _1799_;
assign _1804_ = _1801_ | _1803_;
assign _1805_ = X[156] ^ Y[156];
assign _1806_ = X[156] & Y[156];
assign S[156] = _1805_ ^ _1804_;
assign _1808_ = _1805_ & _1804_;
assign _1809_ = _1806_ | _1808_;
assign _1810_ = X[157] ^ Y[157];
assign _1811_ = X[157] & Y[157];
assign S[157] = _1810_ ^ _1809_;
assign _1813_ = _1810_ & _1809_;
assign _1814_ = _1811_ | _1813_;
assign _1815_ = X[158] ^ Y[158];
assign _1816_ = X[158] & Y[158];
assign S[158] = _1815_ ^ _1814_;
assign _1818_ = _1815_ & _1814_;
assign _1819_ = _1816_ | _1818_;
assign _1820_ = X[159] ^ Y[159];
assign _1821_ = X[159] & Y[159];
assign S[159] = _1820_ ^ _1819_;
assign _1823_ = _1820_ & _1819_;
assign _1824_ = _1821_ | _1823_;
assign _1825_ = X[160] ^ Y[160];
assign _1826_ = X[160] & Y[160];
assign S[160] = _1825_ ^ _1824_;
assign _1828_ = _1825_ & _1824_;
assign _1829_ = _1826_ | _1828_;
assign _1830_ = X[161] ^ Y[161];
assign _1831_ = X[161] & Y[161];
assign S[161] = _1830_ ^ _1829_;
assign _1833_ = _1830_ & _1829_;
assign _1834_ = _1831_ | _1833_;
assign _1835_ = X[162] ^ Y[162];
assign _1836_ = X[162] & Y[162];
assign S[162] = _1835_ ^ _1834_;
assign _1838_ = _1835_ & _1834_;
assign _1839_ = _1836_ | _1838_;
assign _1840_ = X[163] ^ Y[163];
assign _1841_ = X[163] & Y[163];
assign S[163] = _1840_ ^ _1839_;
assign _1843_ = _1840_ & _1839_;
assign _1844_ = _1841_ | _1843_;
assign _1845_ = X[164] ^ Y[164];
assign _1846_ = X[164] & Y[164];
assign S[164] = _1845_ ^ _1844_;
assign _1848_ = _1845_ & _1844_;
assign _1849_ = _1846_ | _1848_;
assign _1850_ = X[165] ^ Y[165];
assign _1851_ = X[165] & Y[165];
assign S[165] = _1850_ ^ _1849_;
assign _1853_ = _1850_ & _1849_;
assign _1854_ = _1851_ | _1853_;
assign _1855_ = X[166] ^ Y[166];
assign _1856_ = X[166] & Y[166];
assign S[166] = _1855_ ^ _1854_;
assign _1858_ = _1855_ & _1854_;
assign _1859_ = _1856_ | _1858_;
assign _1860_ = X[167] ^ Y[167];
assign _1861_ = X[167] & Y[167];
assign S[167] = _1860_ ^ _1859_;
assign _1863_ = _1860_ & _1859_;
assign _1864_ = _1861_ | _1863_;
assign _1865_ = X[168] ^ Y[168];
assign _1866_ = X[168] & Y[168];
assign S[168] = _1865_ ^ _1864_;
assign _1868_ = _1865_ & _1864_;
assign _1869_ = _1866_ | _1868_;
assign _1870_ = X[169] ^ Y[169];
assign _1871_ = X[169] & Y[169];
assign S[169] = _1870_ ^ _1869_;
assign _1873_ = _1870_ & _1869_;
assign _1874_ = _1871_ | _1873_;
assign _1875_ = X[170] ^ Y[170];
assign _1876_ = X[170] & Y[170];
assign S[170] = _1875_ ^ _1874_;
assign _1878_ = _1875_ & _1874_;
assign _1879_ = _1876_ | _1878_;
assign _1880_ = X[171] ^ Y[171];
assign _1881_ = X[171] & Y[171];
assign S[171] = _1880_ ^ _1879_;
assign _1883_ = _1880_ & _1879_;
assign _1884_ = _1881_ | _1883_;
assign _1885_ = X[172] ^ Y[172];
assign _1886_ = X[172] & Y[172];
assign S[172] = _1885_ ^ _1884_;
assign _1888_ = _1885_ & _1884_;
assign _1889_ = _1886_ | _1888_;
assign _1890_ = X[173] ^ Y[173];
assign _1891_ = X[173] & Y[173];
assign S[173] = _1890_ ^ _1889_;
assign _1893_ = _1890_ & _1889_;
assign _1894_ = _1891_ | _1893_;
assign _1895_ = X[174] ^ Y[174];
assign _1896_ = X[174] & Y[174];
assign S[174] = _1895_ ^ _1894_;
assign _1898_ = _1895_ & _1894_;
assign _1899_ = _1896_ | _1898_;
assign _1900_ = X[175] ^ Y[175];
assign _1901_ = X[175] & Y[175];
assign S[175] = _1900_ ^ _1899_;
assign _1903_ = _1900_ & _1899_;
assign _1904_ = _1901_ | _1903_;
assign _1905_ = X[176] ^ Y[176];
assign _1906_ = X[176] & Y[176];
assign S[176] = _1905_ ^ _1904_;
assign _1908_ = _1905_ & _1904_;
assign _1909_ = _1906_ | _1908_;
assign _1910_ = X[177] ^ Y[177];
assign _1911_ = X[177] & Y[177];
assign S[177] = _1910_ ^ _1909_;
assign _1913_ = _1910_ & _1909_;
assign _1914_ = _1911_ | _1913_;
assign _1915_ = X[178] ^ Y[178];
assign _1916_ = X[178] & Y[178];
assign S[178] = _1915_ ^ _1914_;
assign _1918_ = _1915_ & _1914_;
assign _1919_ = _1916_ | _1918_;
assign _1920_ = X[179] ^ Y[179];
assign _1921_ = X[179] & Y[179];
assign S[179] = _1920_ ^ _1919_;
assign _1923_ = _1920_ & _1919_;
assign _1924_ = _1921_ | _1923_;
assign _1925_ = X[180] ^ Y[180];
assign _1926_ = X[180] & Y[180];
assign S[180] = _1925_ ^ _1924_;
assign _1928_ = _1925_ & _1924_;
assign _1929_ = _1926_ | _1928_;
assign _1930_ = X[181] ^ Y[181];
assign _1931_ = X[181] & Y[181];
assign S[181] = _1930_ ^ _1929_;
assign _1933_ = _1930_ & _1929_;
assign _1934_ = _1931_ | _1933_;
assign _1935_ = X[182] ^ Y[182];
assign _1936_ = X[182] & Y[182];
assign S[182] = _1935_ ^ _1934_;
assign _1938_ = _1935_ & _1934_;
assign _1939_ = _1936_ | _1938_;
assign _1940_ = X[183] ^ Y[183];
assign _1941_ = X[183] & Y[183];
assign S[183] = _1940_ ^ _1939_;
assign _1943_ = _1940_ & _1939_;
assign _1944_ = _1941_ | _1943_;
assign _1945_ = X[184] ^ Y[184];
assign _1946_ = X[184] & Y[184];
assign S[184] = _1945_ ^ _1944_;
assign _1948_ = _1945_ & _1944_;
assign _1949_ = _1946_ | _1948_;
assign _1950_ = X[185] ^ Y[185];
assign _1951_ = X[185] & Y[185];
assign S[185] = _1950_ ^ _1949_;
assign _1953_ = _1950_ & _1949_;
assign _1954_ = _1951_ | _1953_;
assign _1955_ = X[186] ^ Y[186];
assign _1956_ = X[186] & Y[186];
assign S[186] = _1955_ ^ _1954_;
assign _1958_ = _1955_ & _1954_;
assign _1959_ = _1956_ | _1958_;
assign _1960_ = X[187] ^ Y[187];
assign _1961_ = X[187] & Y[187];
assign S[187] = _1960_ ^ _1959_;
assign _1963_ = _1960_ & _1959_;
assign _1964_ = _1961_ | _1963_;
assign _1965_ = X[188] ^ Y[188];
assign _1966_ = X[188] & Y[188];
assign S[188] = _1965_ ^ _1964_;
assign _1968_ = _1965_ & _1964_;
assign _1969_ = _1966_ | _1968_;
assign _1970_ = X[189] ^ Y[189];
assign _1971_ = X[189] & Y[189];
assign S[189] = _1970_ ^ _1969_;
assign _1973_ = _1970_ & _1969_;
assign _1974_ = _1971_ | _1973_;
assign _1975_ = X[190] ^ Y[190];
assign _1976_ = X[190] & Y[190];
assign S[190] = _1975_ ^ _1974_;
assign _1978_ = _1975_ & _1974_;
assign _1979_ = _1976_ | _1978_;
assign _1980_ = X[191] ^ Y[191];
assign _1981_ = X[191] & Y[191];
assign S[191] = _1980_ ^ _1979_;
assign _1983_ = _1980_ & _1979_;
assign _1984_ = _1981_ | _1983_;
assign _1985_ = X[192] ^ Y[192];
assign _1986_ = X[192] & Y[192];
assign S[192] = _1985_ ^ _1984_;
assign _1988_ = _1985_ & _1984_;
assign _1989_ = _1986_ | _1988_;
assign _1990_ = X[193] ^ Y[193];
assign _1991_ = X[193] & Y[193];
assign S[193] = _1990_ ^ _1989_;
assign _1993_ = _1990_ & _1989_;
assign _1994_ = _1991_ | _1993_;
assign _1995_ = X[194] ^ Y[194];
assign _1996_ = X[194] & Y[194];
assign S[194] = _1995_ ^ _1994_;
assign _1998_ = _1995_ & _1994_;
assign _1999_ = _1996_ | _1998_;
assign _2000_ = X[195] ^ Y[195];
assign _2001_ = X[195] & Y[195];
assign S[195] = _2000_ ^ _1999_;
assign _2003_ = _2000_ & _1999_;
assign _2004_ = _2001_ | _2003_;
assign _2005_ = X[196] ^ Y[196];
assign _2006_ = X[196] & Y[196];
assign S[196] = _2005_ ^ _2004_;
assign _2008_ = _2005_ & _2004_;
assign _2009_ = _2006_ | _2008_;
assign _2010_ = X[197] ^ Y[197];
assign _2011_ = X[197] & Y[197];
assign S[197] = _2010_ ^ _2009_;
assign _2013_ = _2010_ & _2009_;
assign _2014_ = _2011_ | _2013_;
assign _2015_ = X[198] ^ Y[198];
assign _2016_ = X[198] & Y[198];
assign S[198] = _2015_ ^ _2014_;
assign _2018_ = _2015_ & _2014_;
assign _2019_ = _2016_ | _2018_;
assign _2020_ = X[199] ^ Y[199];
assign _2021_ = X[199] & Y[199];
assign S[199] = _2020_ ^ _2019_;
assign _2023_ = _2020_ & _2019_;
assign _2024_ = _2021_ | _2023_;
assign _2025_ = X[200] ^ Y[200];
assign _2026_ = X[200] & Y[200];
assign S[200] = _2025_ ^ _2024_;
assign _2028_ = _2025_ & _2024_;
assign _2029_ = _2026_ | _2028_;
assign _2030_ = X[201] ^ Y[201];
assign _2031_ = X[201] & Y[201];
assign S[201] = _2030_ ^ _2029_;
assign _2033_ = _2030_ & _2029_;
assign _2034_ = _2031_ | _2033_;
assign _2035_ = X[202] ^ Y[202];
assign _2036_ = X[202] & Y[202];
assign S[202] = _2035_ ^ _2034_;
assign _2038_ = _2035_ & _2034_;
assign _2039_ = _2036_ | _2038_;
assign _2040_ = X[203] ^ Y[203];
assign _2041_ = X[203] & Y[203];
assign S[203] = _2040_ ^ _2039_;
assign _2043_ = _2040_ & _2039_;
assign _2044_ = _2041_ | _2043_;
assign _2045_ = X[204] ^ Y[204];
assign _2046_ = X[204] & Y[204];
assign S[204] = _2045_ ^ _2044_;
assign _2048_ = _2045_ & _2044_;
assign _2049_ = _2046_ | _2048_;
assign _2050_ = X[205] ^ Y[205];
assign _2051_ = X[205] & Y[205];
assign S[205] = _2050_ ^ _2049_;
assign _2053_ = _2050_ & _2049_;
assign _2054_ = _2051_ | _2053_;
assign _2055_ = X[206] ^ Y[206];
assign _2056_ = X[206] & Y[206];
assign S[206] = _2055_ ^ _2054_;
assign _2058_ = _2055_ & _2054_;
assign _2059_ = _2056_ | _2058_;
assign _2060_ = X[207] ^ Y[207];
assign _2061_ = X[207] & Y[207];
assign S[207] = _2060_ ^ _2059_;
assign _2063_ = _2060_ & _2059_;
assign _2064_ = _2061_ | _2063_;
assign _2065_ = X[208] ^ Y[208];
assign _2066_ = X[208] & Y[208];
assign S[208] = _2065_ ^ _2064_;
assign _2068_ = _2065_ & _2064_;
assign _2069_ = _2066_ | _2068_;
assign _2070_ = X[209] ^ Y[209];
assign _2071_ = X[209] & Y[209];
assign S[209] = _2070_ ^ _2069_;
assign _2073_ = _2070_ & _2069_;
assign _2074_ = _2071_ | _2073_;
assign _2075_ = X[210] ^ Y[210];
assign _2076_ = X[210] & Y[210];
assign S[210] = _2075_ ^ _2074_;
assign _2078_ = _2075_ & _2074_;
assign _2079_ = _2076_ | _2078_;
assign _2080_ = X[211] ^ Y[211];
assign _2081_ = X[211] & Y[211];
assign S[211] = _2080_ ^ _2079_;
assign _2083_ = _2080_ & _2079_;
assign _2084_ = _2081_ | _2083_;
assign _2085_ = X[212] ^ Y[212];
assign _2086_ = X[212] & Y[212];
assign S[212] = _2085_ ^ _2084_;
assign _2088_ = _2085_ & _2084_;
assign _2089_ = _2086_ | _2088_;
assign _2090_ = X[213] ^ Y[213];
assign _2091_ = X[213] & Y[213];
assign S[213] = _2090_ ^ _2089_;
assign _2093_ = _2090_ & _2089_;
assign _2094_ = _2091_ | _2093_;
assign _2095_ = X[214] ^ Y[214];
assign _2096_ = X[214] & Y[214];
assign S[214] = _2095_ ^ _2094_;
assign _2098_ = _2095_ & _2094_;
assign _2099_ = _2096_ | _2098_;
assign _2100_ = X[215] ^ Y[215];
assign _2101_ = X[215] & Y[215];
assign S[215] = _2100_ ^ _2099_;
assign _2103_ = _2100_ & _2099_;
assign _2104_ = _2101_ | _2103_;
assign _2105_ = X[216] ^ Y[216];
assign _2106_ = X[216] & Y[216];
assign S[216] = _2105_ ^ _2104_;
assign _2108_ = _2105_ & _2104_;
assign _2109_ = _2106_ | _2108_;
assign _2110_ = X[217] ^ Y[217];
assign _2111_ = X[217] & Y[217];
assign S[217] = _2110_ ^ _2109_;
assign _2113_ = _2110_ & _2109_;
assign _2114_ = _2111_ | _2113_;
assign _2115_ = X[218] ^ Y[218];
assign _2116_ = X[218] & Y[218];
assign S[218] = _2115_ ^ _2114_;
assign _2118_ = _2115_ & _2114_;
assign _2119_ = _2116_ | _2118_;
assign _2120_ = X[219] ^ Y[219];
assign _2121_ = X[219] & Y[219];
assign S[219] = _2120_ ^ _2119_;
assign _2123_ = _2120_ & _2119_;
assign _2124_ = _2121_ | _2123_;
assign _2125_ = X[220] ^ Y[220];
assign _2126_ = X[220] & Y[220];
assign S[220] = _2125_ ^ _2124_;
assign _2128_ = _2125_ & _2124_;
assign _2129_ = _2126_ | _2128_;
assign _2130_ = X[221] ^ Y[221];
assign _2131_ = X[221] & Y[221];
assign S[221] = _2130_ ^ _2129_;
assign _2133_ = _2130_ & _2129_;
assign _2134_ = _2131_ | _2133_;
assign _2135_ = X[222] ^ Y[222];
assign _2136_ = X[222] & Y[222];
assign S[222] = _2135_ ^ _2134_;
assign _2138_ = _2135_ & _2134_;
assign _2139_ = _2136_ | _2138_;
assign _2140_ = X[223] ^ Y[223];
assign _2141_ = X[223] & Y[223];
assign S[223] = _2140_ ^ _2139_;
assign _2143_ = _2140_ & _2139_;
assign _2144_ = _2141_ | _2143_;
assign _2145_ = X[224] ^ Y[224];
assign _2146_ = X[224] & Y[224];
assign S[224] = _2145_ ^ _2144_;
assign _2148_ = _2145_ & _2144_;
assign _2149_ = _2146_ | _2148_;
assign _2150_ = X[225] ^ Y[225];
assign _2151_ = X[225] & Y[225];
assign S[225] = _2150_ ^ _2149_;
assign _2153_ = _2150_ & _2149_;
assign _2154_ = _2151_ | _2153_;
assign _2155_ = X[226] ^ Y[226];
assign _2156_ = X[226] & Y[226];
assign S[226] = _2155_ ^ _2154_;
assign _2158_ = _2155_ & _2154_;
assign _2159_ = _2156_ | _2158_;
assign _2160_ = X[227] ^ Y[227];
assign _2161_ = X[227] & Y[227];
assign S[227] = _2160_ ^ _2159_;
assign _2163_ = _2160_ & _2159_;
assign _2164_ = _2161_ | _2163_;
assign _2165_ = X[228] ^ Y[228];
assign _2166_ = X[228] & Y[228];
assign S[228] = _2165_ ^ _2164_;
assign _2168_ = _2165_ & _2164_;
assign _2169_ = _2166_ | _2168_;
assign _2170_ = X[229] ^ Y[229];
assign _2171_ = X[229] & Y[229];
assign S[229] = _2170_ ^ _2169_;
assign _2173_ = _2170_ & _2169_;
assign _2174_ = _2171_ | _2173_;
assign _2175_ = X[230] ^ Y[230];
assign _2176_ = X[230] & Y[230];
assign S[230] = _2175_ ^ _2174_;
assign _2178_ = _2175_ & _2174_;
assign _2179_ = _2176_ | _2178_;
assign _2180_ = X[231] ^ Y[231];
assign _2181_ = X[231] & Y[231];
assign S[231] = _2180_ ^ _2179_;
assign _2183_ = _2180_ & _2179_;
assign _2184_ = _2181_ | _2183_;
assign _2185_ = X[232] ^ Y[232];
assign _2186_ = X[232] & Y[232];
assign S[232] = _2185_ ^ _2184_;
assign _2188_ = _2185_ & _2184_;
assign _2189_ = _2186_ | _2188_;
assign _2190_ = X[233] ^ Y[233];
assign _2191_ = X[233] & Y[233];
assign S[233] = _2190_ ^ _2189_;
assign _2193_ = _2190_ & _2189_;
assign _2194_ = _2191_ | _2193_;
assign _2195_ = X[234] ^ Y[234];
assign _2196_ = X[234] & Y[234];
assign S[234] = _2195_ ^ _2194_;
assign _2198_ = _2195_ & _2194_;
assign _2199_ = _2196_ | _2198_;
assign _2200_ = X[235] ^ Y[235];
assign _2201_ = X[235] & Y[235];
assign S[235] = _2200_ ^ _2199_;
assign _2203_ = _2200_ & _2199_;
assign _2204_ = _2201_ | _2203_;
assign _2205_ = X[236] ^ Y[236];
assign _2206_ = X[236] & Y[236];
assign S[236] = _2205_ ^ _2204_;
assign _2208_ = _2205_ & _2204_;
assign _2209_ = _2206_ | _2208_;
assign _2210_ = X[237] ^ Y[237];
assign _2211_ = X[237] & Y[237];
assign S[237] = _2210_ ^ _2209_;
assign _2213_ = _2210_ & _2209_;
assign _2214_ = _2211_ | _2213_;
assign _2215_ = X[238] ^ Y[238];
assign _2216_ = X[238] & Y[238];
assign S[238] = _2215_ ^ _2214_;
assign _2218_ = _2215_ & _2214_;
assign _2219_ = _2216_ | _2218_;
assign _2220_ = X[239] ^ Y[239];
assign _2221_ = X[239] & Y[239];
assign S[239] = _2220_ ^ _2219_;
assign _2223_ = _2220_ & _2219_;
assign _2224_ = _2221_ | _2223_;
assign _2225_ = X[240] ^ Y[240];
assign _2226_ = X[240] & Y[240];
assign S[240] = _2225_ ^ _2224_;
assign _2228_ = _2225_ & _2224_;
assign _2229_ = _2226_ | _2228_;
assign _2230_ = X[241] ^ Y[241];
assign _2231_ = X[241] & Y[241];
assign S[241] = _2230_ ^ _2229_;
assign _2233_ = _2230_ & _2229_;
assign _2234_ = _2231_ | _2233_;
assign _2235_ = X[242] ^ Y[242];
assign _2236_ = X[242] & Y[242];
assign S[242] = _2235_ ^ _2234_;
assign _2238_ = _2235_ & _2234_;
assign _2239_ = _2236_ | _2238_;
assign _2240_ = X[243] ^ Y[243];
assign _2241_ = X[243] & Y[243];
assign S[243] = _2240_ ^ _2239_;
assign _2243_ = _2240_ & _2239_;
assign _2244_ = _2241_ | _2243_;
assign _2245_ = X[244] ^ Y[244];
assign _2246_ = X[244] & Y[244];
assign S[244] = _2245_ ^ _2244_;
assign _2248_ = _2245_ & _2244_;
assign _2249_ = _2246_ | _2248_;
assign _2250_ = X[245] ^ Y[245];
assign _2251_ = X[245] & Y[245];
assign S[245] = _2250_ ^ _2249_;
assign _2253_ = _2250_ & _2249_;
assign _2254_ = _2251_ | _2253_;
assign _2255_ = X[246] ^ Y[246];
assign _2256_ = X[246] & Y[246];
assign S[246] = _2255_ ^ _2254_;
assign _2258_ = _2255_ & _2254_;
assign _2259_ = _2256_ | _2258_;
assign _2260_ = X[247] ^ Y[247];
assign _2261_ = X[247] & Y[247];
assign S[247] = _2260_ ^ _2259_;
assign _2263_ = _2260_ & _2259_;
assign _2264_ = _2261_ | _2263_;
assign _2265_ = X[248] ^ Y[248];
assign _2266_ = X[248] & Y[248];
assign S[248] = _2265_ ^ _2264_;
assign _2268_ = _2265_ & _2264_;
assign _2269_ = _2266_ | _2268_;
assign _2270_ = X[249] ^ Y[249];
assign _2271_ = X[249] & Y[249];
assign S[249] = _2270_ ^ _2269_;
assign _2273_ = _2270_ & _2269_;
assign _2274_ = _2271_ | _2273_;
assign _2275_ = X[250] ^ Y[250];
assign _2276_ = X[250] & Y[250];
assign S[250] = _2275_ ^ _2274_;
assign _2278_ = _2275_ & _2274_;
assign _2279_ = _2276_ | _2278_;
assign _2280_ = X[251] ^ Y[251];
assign _2281_ = X[251] & Y[251];
assign S[251] = _2280_ ^ _2279_;
assign _2283_ = _2280_ & _2279_;
assign _2284_ = _2281_ | _2283_;
assign _2285_ = X[252] ^ Y[252];
assign _2286_ = X[252] & Y[252];
assign S[252] = _2285_ ^ _2284_;
assign _2288_ = _2285_ & _2284_;
assign _2289_ = _2286_ | _2288_;
assign _2290_ = X[253] ^ Y[253];
assign _2291_ = X[253] & Y[253];
assign S[253] = _2290_ ^ _2289_;
assign _2293_ = _2290_ & _2289_;
assign _2294_ = _2291_ | _2293_;
assign _2295_ = X[254] ^ Y[254];
assign _2296_ = X[254] & Y[254];
assign S[254] = _2295_ ^ _2294_;
assign _2298_ = _2295_ & _2294_;
assign _2299_ = _2296_ | _2298_;
assign _2300_ = X[255] ^ Y[255];
assign _2301_ = X[255] & Y[255];
assign S[255] = _2300_ ^ _2299_;
assign _2303_ = _2300_ & _2299_;
assign _2304_ = _2301_ | _2303_;
assign _2305_ = X[256] ^ Y[256];
assign _2306_ = X[256] & Y[256];
assign S[256] = _2305_ ^ _2304_;
assign _2308_ = _2305_ & _2304_;
assign _2309_ = _2306_ | _2308_;
assign _2310_ = X[257] ^ Y[257];
assign _2311_ = X[257] & Y[257];
assign S[257] = _2310_ ^ _2309_;
assign _2313_ = _2310_ & _2309_;
assign _2314_ = _2311_ | _2313_;
assign _2315_ = X[258] ^ Y[258];
assign _2316_ = X[258] & Y[258];
assign S[258] = _2315_ ^ _2314_;
assign _2318_ = _2315_ & _2314_;
assign _2319_ = _2316_ | _2318_;
assign _2320_ = X[259] ^ Y[259];
assign _2321_ = X[259] & Y[259];
assign S[259] = _2320_ ^ _2319_;
assign _2323_ = _2320_ & _2319_;
assign _2324_ = _2321_ | _2323_;
assign _2325_ = X[260] ^ Y[260];
assign _2326_ = X[260] & Y[260];
assign S[260] = _2325_ ^ _2324_;
assign _2328_ = _2325_ & _2324_;
assign _2329_ = _2326_ | _2328_;
assign _2330_ = X[261] ^ Y[261];
assign _2331_ = X[261] & Y[261];
assign S[261] = _2330_ ^ _2329_;
assign _2333_ = _2330_ & _2329_;
assign _2334_ = _2331_ | _2333_;
assign _2335_ = X[262] ^ Y[262];
assign _2336_ = X[262] & Y[262];
assign S[262] = _2335_ ^ _2334_;
assign _2338_ = _2335_ & _2334_;
assign _2339_ = _2336_ | _2338_;
assign _2340_ = X[263] ^ Y[263];
assign _2341_ = X[263] & Y[263];
assign S[263] = _2340_ ^ _2339_;
assign _2343_ = _2340_ & _2339_;
assign _2344_ = _2341_ | _2343_;
assign _2345_ = X[264] ^ Y[264];
assign _2346_ = X[264] & Y[264];
assign S[264] = _2345_ ^ _2344_;
assign _2348_ = _2345_ & _2344_;
assign _2349_ = _2346_ | _2348_;
assign _2350_ = X[265] ^ Y[265];
assign _2351_ = X[265] & Y[265];
assign S[265] = _2350_ ^ _2349_;
assign _2353_ = _2350_ & _2349_;
assign _2354_ = _2351_ | _2353_;
assign _2355_ = X[266] ^ Y[266];
assign _2356_ = X[266] & Y[266];
assign S[266] = _2355_ ^ _2354_;
assign _2358_ = _2355_ & _2354_;
assign _2359_ = _2356_ | _2358_;
assign _2360_ = X[267] ^ Y[267];
assign _2361_ = X[267] & Y[267];
assign S[267] = _2360_ ^ _2359_;
assign _2363_ = _2360_ & _2359_;
assign _2364_ = _2361_ | _2363_;
assign _2365_ = X[268] ^ Y[268];
assign _2366_ = X[268] & Y[268];
assign S[268] = _2365_ ^ _2364_;
assign _2368_ = _2365_ & _2364_;
assign _2369_ = _2366_ | _2368_;
assign _2370_ = X[269] ^ Y[269];
assign _2371_ = X[269] & Y[269];
assign S[269] = _2370_ ^ _2369_;
assign _2373_ = _2370_ & _2369_;
assign _2374_ = _2371_ | _2373_;
assign _2375_ = X[270] ^ Y[270];
assign _2376_ = X[270] & Y[270];
assign S[270] = _2375_ ^ _2374_;
assign _2378_ = _2375_ & _2374_;
assign _2379_ = _2376_ | _2378_;
assign _2380_ = X[271] ^ Y[271];
assign _2381_ = X[271] & Y[271];
assign S[271] = _2380_ ^ _2379_;
assign _2383_ = _2380_ & _2379_;
assign _2384_ = _2381_ | _2383_;
assign _2385_ = X[272] ^ Y[272];
assign _2386_ = X[272] & Y[272];
assign S[272] = _2385_ ^ _2384_;
assign _2388_ = _2385_ & _2384_;
assign _2389_ = _2386_ | _2388_;
assign _2390_ = X[273] ^ Y[273];
assign _2391_ = X[273] & Y[273];
assign S[273] = _2390_ ^ _2389_;
assign _2393_ = _2390_ & _2389_;
assign _2394_ = _2391_ | _2393_;
assign _2395_ = X[274] ^ Y[274];
assign _2396_ = X[274] & Y[274];
assign S[274] = _2395_ ^ _2394_;
assign _2398_ = _2395_ & _2394_;
assign _2399_ = _2396_ | _2398_;
assign _2400_ = X[275] ^ Y[275];
assign _2401_ = X[275] & Y[275];
assign S[275] = _2400_ ^ _2399_;
assign _2403_ = _2400_ & _2399_;
assign _2404_ = _2401_ | _2403_;
assign _2405_ = X[276] ^ Y[276];
assign _2406_ = X[276] & Y[276];
assign S[276] = _2405_ ^ _2404_;
assign _2408_ = _2405_ & _2404_;
assign _2409_ = _2406_ | _2408_;
assign _2410_ = X[277] ^ Y[277];
assign _2411_ = X[277] & Y[277];
assign S[277] = _2410_ ^ _2409_;
assign _2413_ = _2410_ & _2409_;
assign _2414_ = _2411_ | _2413_;
assign _2415_ = X[278] ^ Y[278];
assign _2416_ = X[278] & Y[278];
assign S[278] = _2415_ ^ _2414_;
assign _2418_ = _2415_ & _2414_;
assign _2419_ = _2416_ | _2418_;
assign _2420_ = X[279] ^ Y[279];
assign _2421_ = X[279] & Y[279];
assign S[279] = _2420_ ^ _2419_;
assign _2423_ = _2420_ & _2419_;
assign _2424_ = _2421_ | _2423_;
assign _2425_ = X[280] ^ Y[280];
assign _2426_ = X[280] & Y[280];
assign S[280] = _2425_ ^ _2424_;
assign _2428_ = _2425_ & _2424_;
assign _2429_ = _2426_ | _2428_;
assign _2430_ = X[281] ^ Y[281];
assign _2431_ = X[281] & Y[281];
assign S[281] = _2430_ ^ _2429_;
assign _2433_ = _2430_ & _2429_;
assign _2434_ = _2431_ | _2433_;
assign _2435_ = X[282] ^ Y[282];
assign _2436_ = X[282] & Y[282];
assign S[282] = _2435_ ^ _2434_;
assign _2438_ = _2435_ & _2434_;
assign _2439_ = _2436_ | _2438_;
assign _2440_ = X[283] ^ Y[283];
assign _2441_ = X[283] & Y[283];
assign S[283] = _2440_ ^ _2439_;
assign _2443_ = _2440_ & _2439_;
assign _2444_ = _2441_ | _2443_;
assign _2445_ = X[284] ^ Y[284];
assign _2446_ = X[284] & Y[284];
assign S[284] = _2445_ ^ _2444_;
assign _2448_ = _2445_ & _2444_;
assign _2449_ = _2446_ | _2448_;
assign _2450_ = X[285] ^ Y[285];
assign _2451_ = X[285] & Y[285];
assign S[285] = _2450_ ^ _2449_;
assign _2453_ = _2450_ & _2449_;
assign _2454_ = _2451_ | _2453_;
assign _2455_ = X[286] ^ Y[286];
assign _2456_ = X[286] & Y[286];
assign S[286] = _2455_ ^ _2454_;
assign _2458_ = _2455_ & _2454_;
assign _2459_ = _2456_ | _2458_;
assign _2460_ = X[287] ^ Y[287];
assign _2461_ = X[287] & Y[287];
assign S[287] = _2460_ ^ _2459_;
assign _2463_ = _2460_ & _2459_;
assign _2464_ = _2461_ | _2463_;
assign _2465_ = X[288] ^ Y[288];
assign _2466_ = X[288] & Y[288];
assign S[288] = _2465_ ^ _2464_;
assign _2468_ = _2465_ & _2464_;
assign _2469_ = _2466_ | _2468_;
assign _2470_ = X[289] ^ Y[289];
assign _2471_ = X[289] & Y[289];
assign S[289] = _2470_ ^ _2469_;
assign _2473_ = _2470_ & _2469_;
assign _2474_ = _2471_ | _2473_;
assign _2475_ = X[290] ^ Y[290];
assign _2476_ = X[290] & Y[290];
assign S[290] = _2475_ ^ _2474_;
assign _2478_ = _2475_ & _2474_;
assign _2479_ = _2476_ | _2478_;
assign _2480_ = X[291] ^ Y[291];
assign _2481_ = X[291] & Y[291];
assign S[291] = _2480_ ^ _2479_;
assign _2483_ = _2480_ & _2479_;
assign _2484_ = _2481_ | _2483_;
assign _2485_ = X[292] ^ Y[292];
assign _2486_ = X[292] & Y[292];
assign S[292] = _2485_ ^ _2484_;
assign _2488_ = _2485_ & _2484_;
assign _2489_ = _2486_ | _2488_;
assign _2490_ = X[293] ^ Y[293];
assign _2491_ = X[293] & Y[293];
assign S[293] = _2490_ ^ _2489_;
assign _2493_ = _2490_ & _2489_;
assign _2494_ = _2491_ | _2493_;
assign _2495_ = X[294] ^ Y[294];
assign _2496_ = X[294] & Y[294];
assign S[294] = _2495_ ^ _2494_;
assign _2498_ = _2495_ & _2494_;
assign _2499_ = _2496_ | _2498_;
assign _2500_ = X[295] ^ Y[295];
assign _2501_ = X[295] & Y[295];
assign S[295] = _2500_ ^ _2499_;
assign _2503_ = _2500_ & _2499_;
assign _2504_ = _2501_ | _2503_;
assign _2505_ = X[296] ^ Y[296];
assign _2506_ = X[296] & Y[296];
assign S[296] = _2505_ ^ _2504_;
assign _2508_ = _2505_ & _2504_;
assign _2509_ = _2506_ | _2508_;
assign _2510_ = X[297] ^ Y[297];
assign _2511_ = X[297] & Y[297];
assign S[297] = _2510_ ^ _2509_;
assign _2513_ = _2510_ & _2509_;
assign _2514_ = _2511_ | _2513_;
assign _2515_ = X[298] ^ Y[298];
assign _2516_ = X[298] & Y[298];
assign S[298] = _2515_ ^ _2514_;
assign _2518_ = _2515_ & _2514_;
assign _2519_ = _2516_ | _2518_;
assign _2520_ = X[299] ^ Y[299];
assign _2521_ = X[299] & Y[299];
assign S[299] = _2520_ ^ _2519_;
assign _2523_ = _2520_ & _2519_;
assign _2524_ = _2521_ | _2523_;
assign _2525_ = X[300] ^ Y[300];
assign _2526_ = X[300] & Y[300];
assign S[300] = _2525_ ^ _2524_;
assign _2528_ = _2525_ & _2524_;
assign _2529_ = _2526_ | _2528_;
assign _2530_ = X[301] ^ Y[301];
assign _2531_ = X[301] & Y[301];
assign S[301] = _2530_ ^ _2529_;
assign _2533_ = _2530_ & _2529_;
assign _2534_ = _2531_ | _2533_;
assign _2535_ = X[302] ^ Y[302];
assign _2536_ = X[302] & Y[302];
assign S[302] = _2535_ ^ _2534_;
assign _2538_ = _2535_ & _2534_;
assign _2539_ = _2536_ | _2538_;
assign _2540_ = X[303] ^ Y[303];
assign _2541_ = X[303] & Y[303];
assign S[303] = _2540_ ^ _2539_;
assign _2543_ = _2540_ & _2539_;
assign _2544_ = _2541_ | _2543_;
assign _2545_ = X[304] ^ Y[304];
assign _2546_ = X[304] & Y[304];
assign S[304] = _2545_ ^ _2544_;
assign _2548_ = _2545_ & _2544_;
assign _2549_ = _2546_ | _2548_;
assign _2550_ = X[305] ^ Y[305];
assign _2551_ = X[305] & Y[305];
assign S[305] = _2550_ ^ _2549_;
assign _2553_ = _2550_ & _2549_;
assign _2554_ = _2551_ | _2553_;
assign _2555_ = X[306] ^ Y[306];
assign _2556_ = X[306] & Y[306];
assign S[306] = _2555_ ^ _2554_;
assign _2558_ = _2555_ & _2554_;
assign _2559_ = _2556_ | _2558_;
assign _2560_ = X[307] ^ Y[307];
assign _2561_ = X[307] & Y[307];
assign S[307] = _2560_ ^ _2559_;
assign _2563_ = _2560_ & _2559_;
assign _2564_ = _2561_ | _2563_;
assign _2565_ = X[308] ^ Y[308];
assign _2566_ = X[308] & Y[308];
assign S[308] = _2565_ ^ _2564_;
assign _2568_ = _2565_ & _2564_;
assign _2569_ = _2566_ | _2568_;
assign _2570_ = X[309] ^ Y[309];
assign _2571_ = X[309] & Y[309];
assign S[309] = _2570_ ^ _2569_;
assign _2573_ = _2570_ & _2569_;
assign _2574_ = _2571_ | _2573_;
assign _2575_ = X[310] ^ Y[310];
assign _2576_ = X[310] & Y[310];
assign S[310] = _2575_ ^ _2574_;
assign _2578_ = _2575_ & _2574_;
assign _2579_ = _2576_ | _2578_;
assign _2580_ = X[311] ^ Y[311];
assign _2581_ = X[311] & Y[311];
assign S[311] = _2580_ ^ _2579_;
assign _2583_ = _2580_ & _2579_;
assign _2584_ = _2581_ | _2583_;
assign _2585_ = X[312] ^ Y[312];
assign _2586_ = X[312] & Y[312];
assign S[312] = _2585_ ^ _2584_;
assign _2588_ = _2585_ & _2584_;
assign _2589_ = _2586_ | _2588_;
assign _2590_ = X[313] ^ Y[313];
assign _2591_ = X[313] & Y[313];
assign S[313] = _2590_ ^ _2589_;
assign _2593_ = _2590_ & _2589_;
assign _2594_ = _2591_ | _2593_;
assign _2595_ = X[314] ^ Y[314];
assign _2596_ = X[314] & Y[314];
assign S[314] = _2595_ ^ _2594_;
assign _2598_ = _2595_ & _2594_;
assign _2599_ = _2596_ | _2598_;
assign _2600_ = X[315] ^ Y[315];
assign _2601_ = X[315] & Y[315];
assign S[315] = _2600_ ^ _2599_;
assign _2603_ = _2600_ & _2599_;
assign _2604_ = _2601_ | _2603_;
assign _2605_ = X[316] ^ Y[316];
assign _2606_ = X[316] & Y[316];
assign S[316] = _2605_ ^ _2604_;
assign _2608_ = _2605_ & _2604_;
assign _2609_ = _2606_ | _2608_;
assign _2610_ = X[317] ^ Y[317];
assign _2611_ = X[317] & Y[317];
assign S[317] = _2610_ ^ _2609_;
assign _2613_ = _2610_ & _2609_;
assign _2614_ = _2611_ | _2613_;
assign _2615_ = X[318] ^ Y[318];
assign _2616_ = X[318] & Y[318];
assign S[318] = _2615_ ^ _2614_;
assign _2618_ = _2615_ & _2614_;
assign _2619_ = _2616_ | _2618_;
assign _2620_ = X[319] ^ Y[319];
assign _2621_ = X[319] & Y[319];
assign S[319] = _2620_ ^ _2619_;
assign _2623_ = _2620_ & _2619_;
assign _2624_ = _2621_ | _2623_;
assign _2625_ = X[320] ^ Y[320];
assign _2626_ = X[320] & Y[320];
assign S[320] = _2625_ ^ _2624_;
assign _2628_ = _2625_ & _2624_;
assign _2629_ = _2626_ | _2628_;
assign _2630_ = X[321] ^ Y[321];
assign _2631_ = X[321] & Y[321];
assign S[321] = _2630_ ^ _2629_;
assign _2633_ = _2630_ & _2629_;
assign _2634_ = _2631_ | _2633_;
assign _2635_ = X[322] ^ Y[322];
assign _2636_ = X[322] & Y[322];
assign S[322] = _2635_ ^ _2634_;
assign _2638_ = _2635_ & _2634_;
assign _2639_ = _2636_ | _2638_;
assign _2640_ = X[323] ^ Y[323];
assign _2641_ = X[323] & Y[323];
assign S[323] = _2640_ ^ _2639_;
assign _2643_ = _2640_ & _2639_;
assign _2644_ = _2641_ | _2643_;
assign _2645_ = X[324] ^ Y[324];
assign _2646_ = X[324] & Y[324];
assign S[324] = _2645_ ^ _2644_;
assign _2648_ = _2645_ & _2644_;
assign _2649_ = _2646_ | _2648_;
assign _2650_ = X[325] ^ Y[325];
assign _2651_ = X[325] & Y[325];
assign S[325] = _2650_ ^ _2649_;
assign _2653_ = _2650_ & _2649_;
assign _2654_ = _2651_ | _2653_;
assign _2655_ = X[326] ^ Y[326];
assign _2656_ = X[326] & Y[326];
assign S[326] = _2655_ ^ _2654_;
assign _2658_ = _2655_ & _2654_;
assign _2659_ = _2656_ | _2658_;
assign _2660_ = X[327] ^ Y[327];
assign _2661_ = X[327] & Y[327];
assign S[327] = _2660_ ^ _2659_;
assign _2663_ = _2660_ & _2659_;
assign _2664_ = _2661_ | _2663_;
assign _2665_ = X[328] ^ Y[328];
assign _2666_ = X[328] & Y[328];
assign S[328] = _2665_ ^ _2664_;
assign _2668_ = _2665_ & _2664_;
assign _2669_ = _2666_ | _2668_;
assign _2670_ = X[329] ^ Y[329];
assign _2671_ = X[329] & Y[329];
assign S[329] = _2670_ ^ _2669_;
assign _2673_ = _2670_ & _2669_;
assign _2674_ = _2671_ | _2673_;
assign _2675_ = X[330] ^ Y[330];
assign _2676_ = X[330] & Y[330];
assign S[330] = _2675_ ^ _2674_;
assign _2678_ = _2675_ & _2674_;
assign _2679_ = _2676_ | _2678_;
assign _2680_ = X[331] ^ Y[331];
assign _2681_ = X[331] & Y[331];
assign S[331] = _2680_ ^ _2679_;
assign _2683_ = _2680_ & _2679_;
assign _2684_ = _2681_ | _2683_;
assign _2685_ = X[332] ^ Y[332];
assign _2686_ = X[332] & Y[332];
assign S[332] = _2685_ ^ _2684_;
assign _2688_ = _2685_ & _2684_;
assign _2689_ = _2686_ | _2688_;
assign _2690_ = X[333] ^ Y[333];
assign _2691_ = X[333] & Y[333];
assign S[333] = _2690_ ^ _2689_;
assign _2693_ = _2690_ & _2689_;
assign _2694_ = _2691_ | _2693_;
assign _2695_ = X[334] ^ Y[334];
assign _2696_ = X[334] & Y[334];
assign S[334] = _2695_ ^ _2694_;
assign _2698_ = _2695_ & _2694_;
assign _2699_ = _2696_ | _2698_;
assign _2700_ = X[335] ^ Y[335];
assign _2701_ = X[335] & Y[335];
assign S[335] = _2700_ ^ _2699_;
assign _2703_ = _2700_ & _2699_;
assign _2704_ = _2701_ | _2703_;
assign _2705_ = X[336] ^ Y[336];
assign _2706_ = X[336] & Y[336];
assign S[336] = _2705_ ^ _2704_;
assign _2708_ = _2705_ & _2704_;
assign _2709_ = _2706_ | _2708_;
assign _2710_ = X[337] ^ Y[337];
assign _2711_ = X[337] & Y[337];
assign S[337] = _2710_ ^ _2709_;
assign _2713_ = _2710_ & _2709_;
assign _2714_ = _2711_ | _2713_;
assign _2715_ = X[338] ^ Y[338];
assign _2716_ = X[338] & Y[338];
assign S[338] = _2715_ ^ _2714_;
assign _2718_ = _2715_ & _2714_;
assign _2719_ = _2716_ | _2718_;
assign _2720_ = X[339] ^ Y[339];
assign _2721_ = X[339] & Y[339];
assign S[339] = _2720_ ^ _2719_;
assign _2723_ = _2720_ & _2719_;
assign _2724_ = _2721_ | _2723_;
assign _2725_ = X[340] ^ Y[340];
assign _2726_ = X[340] & Y[340];
assign S[340] = _2725_ ^ _2724_;
assign _2728_ = _2725_ & _2724_;
assign _2729_ = _2726_ | _2728_;
assign _2730_ = X[341] ^ Y[341];
assign _2731_ = X[341] & Y[341];
assign S[341] = _2730_ ^ _2729_;
assign _2733_ = _2730_ & _2729_;
assign _2734_ = _2731_ | _2733_;
assign _2735_ = X[342] ^ Y[342];
assign _2736_ = X[342] & Y[342];
assign S[342] = _2735_ ^ _2734_;
assign _2738_ = _2735_ & _2734_;
assign _2739_ = _2736_ | _2738_;
assign _2740_ = X[343] ^ Y[343];
assign _2741_ = X[343] & Y[343];
assign S[343] = _2740_ ^ _2739_;
assign _2743_ = _2740_ & _2739_;
assign _2744_ = _2741_ | _2743_;
assign _2745_ = X[344] ^ Y[344];
assign _2746_ = X[344] & Y[344];
assign S[344] = _2745_ ^ _2744_;
assign _2748_ = _2745_ & _2744_;
assign _2749_ = _2746_ | _2748_;
assign _2750_ = X[345] ^ Y[345];
assign _2751_ = X[345] & Y[345];
assign S[345] = _2750_ ^ _2749_;
assign _2753_ = _2750_ & _2749_;
assign _2754_ = _2751_ | _2753_;
assign _2755_ = X[346] ^ Y[346];
assign _2756_ = X[346] & Y[346];
assign S[346] = _2755_ ^ _2754_;
assign _2758_ = _2755_ & _2754_;
assign _2759_ = _2756_ | _2758_;
assign _2760_ = X[347] ^ Y[347];
assign _2761_ = X[347] & Y[347];
assign S[347] = _2760_ ^ _2759_;
assign _2763_ = _2760_ & _2759_;
assign _2764_ = _2761_ | _2763_;
assign _2765_ = X[348] ^ Y[348];
assign _2766_ = X[348] & Y[348];
assign S[348] = _2765_ ^ _2764_;
assign _2768_ = _2765_ & _2764_;
assign _2769_ = _2766_ | _2768_;
assign _2770_ = X[349] ^ Y[349];
assign _2771_ = X[349] & Y[349];
assign S[349] = _2770_ ^ _2769_;
assign _2773_ = _2770_ & _2769_;
assign _2774_ = _2771_ | _2773_;
assign _2775_ = X[350] ^ Y[350];
assign _2776_ = X[350] & Y[350];
assign S[350] = _2775_ ^ _2774_;
assign _2778_ = _2775_ & _2774_;
assign _2779_ = _2776_ | _2778_;
assign _2780_ = X[351] ^ Y[351];
assign _2781_ = X[351] & Y[351];
assign S[351] = _2780_ ^ _2779_;
assign _2783_ = _2780_ & _2779_;
assign _2784_ = _2781_ | _2783_;
assign _2785_ = X[352] ^ Y[352];
assign _2786_ = X[352] & Y[352];
assign S[352] = _2785_ ^ _2784_;
assign _2788_ = _2785_ & _2784_;
assign _2789_ = _2786_ | _2788_;
assign _2790_ = X[353] ^ Y[353];
assign _2791_ = X[353] & Y[353];
assign S[353] = _2790_ ^ _2789_;
assign _2793_ = _2790_ & _2789_;
assign _2794_ = _2791_ | _2793_;
assign _2795_ = X[354] ^ Y[354];
assign _2796_ = X[354] & Y[354];
assign S[354] = _2795_ ^ _2794_;
assign _2798_ = _2795_ & _2794_;
assign _2799_ = _2796_ | _2798_;
assign _2800_ = X[355] ^ Y[355];
assign _2801_ = X[355] & Y[355];
assign S[355] = _2800_ ^ _2799_;
assign _2803_ = _2800_ & _2799_;
assign _2804_ = _2801_ | _2803_;
assign _2805_ = X[356] ^ Y[356];
assign _2806_ = X[356] & Y[356];
assign S[356] = _2805_ ^ _2804_;
assign _2808_ = _2805_ & _2804_;
assign _2809_ = _2806_ | _2808_;
assign _2810_ = X[357] ^ Y[357];
assign _2811_ = X[357] & Y[357];
assign S[357] = _2810_ ^ _2809_;
assign _2813_ = _2810_ & _2809_;
assign _2814_ = _2811_ | _2813_;
assign _2815_ = X[358] ^ Y[358];
assign _2816_ = X[358] & Y[358];
assign S[358] = _2815_ ^ _2814_;
assign _2818_ = _2815_ & _2814_;
assign _2819_ = _2816_ | _2818_;
assign _2820_ = X[359] ^ Y[359];
assign _2821_ = X[359] & Y[359];
assign S[359] = _2820_ ^ _2819_;
assign _2823_ = _2820_ & _2819_;
assign _2824_ = _2821_ | _2823_;
assign _2825_ = X[360] ^ Y[360];
assign _2826_ = X[360] & Y[360];
assign S[360] = _2825_ ^ _2824_;
assign _2828_ = _2825_ & _2824_;
assign _2829_ = _2826_ | _2828_;
assign _2830_ = X[361] ^ Y[361];
assign _2831_ = X[361] & Y[361];
assign S[361] = _2830_ ^ _2829_;
assign _2833_ = _2830_ & _2829_;
assign _2834_ = _2831_ | _2833_;
assign _2835_ = X[362] ^ Y[362];
assign _2836_ = X[362] & Y[362];
assign S[362] = _2835_ ^ _2834_;
assign _2838_ = _2835_ & _2834_;
assign _2839_ = _2836_ | _2838_;
assign _2840_ = X[363] ^ Y[363];
assign _2841_ = X[363] & Y[363];
assign S[363] = _2840_ ^ _2839_;
assign _2843_ = _2840_ & _2839_;
assign _2844_ = _2841_ | _2843_;
assign _2845_ = X[364] ^ Y[364];
assign _2846_ = X[364] & Y[364];
assign S[364] = _2845_ ^ _2844_;
assign _2848_ = _2845_ & _2844_;
assign _2849_ = _2846_ | _2848_;
assign _2850_ = X[365] ^ Y[365];
assign _2851_ = X[365] & Y[365];
assign S[365] = _2850_ ^ _2849_;
assign _2853_ = _2850_ & _2849_;
assign _2854_ = _2851_ | _2853_;
assign _2855_ = X[366] ^ Y[366];
assign _2856_ = X[366] & Y[366];
assign S[366] = _2855_ ^ _2854_;
assign _2858_ = _2855_ & _2854_;
assign _2859_ = _2856_ | _2858_;
assign _2860_ = X[367] ^ Y[367];
assign _2861_ = X[367] & Y[367];
assign S[367] = _2860_ ^ _2859_;
assign _2863_ = _2860_ & _2859_;
assign _2864_ = _2861_ | _2863_;
assign _2865_ = X[368] ^ Y[368];
assign _2866_ = X[368] & Y[368];
assign S[368] = _2865_ ^ _2864_;
assign _2868_ = _2865_ & _2864_;
assign _2869_ = _2866_ | _2868_;
assign _2870_ = X[369] ^ Y[369];
assign _2871_ = X[369] & Y[369];
assign S[369] = _2870_ ^ _2869_;
assign _2873_ = _2870_ & _2869_;
assign _2874_ = _2871_ | _2873_;
assign _2875_ = X[370] ^ Y[370];
assign _2876_ = X[370] & Y[370];
assign S[370] = _2875_ ^ _2874_;
assign _2878_ = _2875_ & _2874_;
assign _2879_ = _2876_ | _2878_;
assign _2880_ = X[371] ^ Y[371];
assign _2881_ = X[371] & Y[371];
assign S[371] = _2880_ ^ _2879_;
assign _2883_ = _2880_ & _2879_;
assign _2884_ = _2881_ | _2883_;
assign _2885_ = X[372] ^ Y[372];
assign _2886_ = X[372] & Y[372];
assign S[372] = _2885_ ^ _2884_;
assign _2888_ = _2885_ & _2884_;
assign _2889_ = _2886_ | _2888_;
assign _2890_ = X[373] ^ Y[373];
assign _2891_ = X[373] & Y[373];
assign S[373] = _2890_ ^ _2889_;
assign _2893_ = _2890_ & _2889_;
assign _2894_ = _2891_ | _2893_;
assign _2895_ = X[374] ^ Y[374];
assign _2896_ = X[374] & Y[374];
assign S[374] = _2895_ ^ _2894_;
assign _2898_ = _2895_ & _2894_;
assign _2899_ = _2896_ | _2898_;
assign _2900_ = X[375] ^ Y[375];
assign _2901_ = X[375] & Y[375];
assign S[375] = _2900_ ^ _2899_;
assign _2903_ = _2900_ & _2899_;
assign _2904_ = _2901_ | _2903_;
assign _2905_ = X[376] ^ Y[376];
assign _2906_ = X[376] & Y[376];
assign S[376] = _2905_ ^ _2904_;
assign _2908_ = _2905_ & _2904_;
assign _2909_ = _2906_ | _2908_;
assign _2910_ = X[377] ^ Y[377];
assign _2911_ = X[377] & Y[377];
assign S[377] = _2910_ ^ _2909_;
assign _2913_ = _2910_ & _2909_;
assign _2914_ = _2911_ | _2913_;
assign _2915_ = X[378] ^ Y[378];
assign _2916_ = X[378] & Y[378];
assign S[378] = _2915_ ^ _2914_;
assign _2918_ = _2915_ & _2914_;
assign _2919_ = _2916_ | _2918_;
assign _2920_ = X[379] ^ Y[379];
assign _2921_ = X[379] & Y[379];
assign S[379] = _2920_ ^ _2919_;
assign _2923_ = _2920_ & _2919_;
assign _2924_ = _2921_ | _2923_;
assign _2925_ = X[380] ^ Y[380];
assign _2926_ = X[380] & Y[380];
assign S[380] = _2925_ ^ _2924_;
assign _2928_ = _2925_ & _2924_;
assign _2929_ = _2926_ | _2928_;
assign _2930_ = X[381] ^ Y[381];
assign _2931_ = X[381] & Y[381];
assign S[381] = _2930_ ^ _2929_;
assign _2933_ = _2930_ & _2929_;
assign _2934_ = _2931_ | _2933_;
assign _2935_ = X[382] ^ Y[382];
assign _2936_ = X[382] & Y[382];
assign S[382] = _2935_ ^ _2934_;
assign _2938_ = _2935_ & _2934_;
assign _2939_ = _2936_ | _2938_;
assign _2940_ = X[383] ^ Y[383];
assign _2941_ = X[383] & Y[383];
assign S[383] = _2940_ ^ _2939_;
assign _2943_ = _2940_ & _2939_;
assign _2944_ = _2941_ | _2943_;
assign _2945_ = X[384] ^ Y[384];
assign _2946_ = X[384] & Y[384];
assign S[384] = _2945_ ^ _2944_;
assign _2948_ = _2945_ & _2944_;
assign _2949_ = _2946_ | _2948_;
assign _2950_ = X[385] ^ Y[385];
assign _2951_ = X[385] & Y[385];
assign S[385] = _2950_ ^ _2949_;
assign _2953_ = _2950_ & _2949_;
assign _2954_ = _2951_ | _2953_;
assign _2955_ = X[386] ^ Y[386];
assign _2956_ = X[386] & Y[386];
assign S[386] = _2955_ ^ _2954_;
assign _2958_ = _2955_ & _2954_;
assign _2959_ = _2956_ | _2958_;
assign _2960_ = X[387] ^ Y[387];
assign _2961_ = X[387] & Y[387];
assign S[387] = _2960_ ^ _2959_;
assign _2963_ = _2960_ & _2959_;
assign _2964_ = _2961_ | _2963_;
assign _2965_ = X[388] ^ Y[388];
assign _2966_ = X[388] & Y[388];
assign S[388] = _2965_ ^ _2964_;
assign _2968_ = _2965_ & _2964_;
assign _2969_ = _2966_ | _2968_;
assign _2970_ = X[389] ^ Y[389];
assign _2971_ = X[389] & Y[389];
assign S[389] = _2970_ ^ _2969_;
assign _2973_ = _2970_ & _2969_;
assign _2974_ = _2971_ | _2973_;
assign _2975_ = X[390] ^ Y[390];
assign _2976_ = X[390] & Y[390];
assign S[390] = _2975_ ^ _2974_;
assign _2978_ = _2975_ & _2974_;
assign _2979_ = _2976_ | _2978_;
assign _2980_ = X[391] ^ Y[391];
assign _2981_ = X[391] & Y[391];
assign S[391] = _2980_ ^ _2979_;
assign _2983_ = _2980_ & _2979_;
assign _2984_ = _2981_ | _2983_;
assign _2985_ = X[392] ^ Y[392];
assign _2986_ = X[392] & Y[392];
assign S[392] = _2985_ ^ _2984_;
assign _2988_ = _2985_ & _2984_;
assign _2989_ = _2986_ | _2988_;
assign _2990_ = X[393] ^ Y[393];
assign _2991_ = X[393] & Y[393];
assign S[393] = _2990_ ^ _2989_;
assign _2993_ = _2990_ & _2989_;
assign _2994_ = _2991_ | _2993_;
assign _2995_ = X[394] ^ Y[394];
assign _2996_ = X[394] & Y[394];
assign S[394] = _2995_ ^ _2994_;
assign _2998_ = _2995_ & _2994_;
assign _2999_ = _2996_ | _2998_;
assign _3000_ = X[395] ^ Y[395];
assign _3001_ = X[395] & Y[395];
assign S[395] = _3000_ ^ _2999_;
assign _3003_ = _3000_ & _2999_;
assign _3004_ = _3001_ | _3003_;
assign _3005_ = X[396] ^ Y[396];
assign _3006_ = X[396] & Y[396];
assign S[396] = _3005_ ^ _3004_;
assign _3008_ = _3005_ & _3004_;
assign _3009_ = _3006_ | _3008_;
assign _3010_ = X[397] ^ Y[397];
assign _3011_ = X[397] & Y[397];
assign S[397] = _3010_ ^ _3009_;
assign _3013_ = _3010_ & _3009_;
assign _3014_ = _3011_ | _3013_;
assign _3015_ = X[398] ^ Y[398];
assign _3016_ = X[398] & Y[398];
assign S[398] = _3015_ ^ _3014_;
assign _3018_ = _3015_ & _3014_;
assign _3019_ = _3016_ | _3018_;
assign _3020_ = X[399] ^ Y[399];
assign _3021_ = X[399] & Y[399];
assign S[399] = _3020_ ^ _3019_;
assign _3023_ = _3020_ & _3019_;
assign _3024_ = _3021_ | _3023_;
assign _3025_ = X[400] ^ Y[400];
assign _3026_ = X[400] & Y[400];
assign S[400] = _3025_ ^ _3024_;
assign _3028_ = _3025_ & _3024_;
assign _3029_ = _3026_ | _3028_;
assign _3030_ = X[401] ^ Y[401];
assign _3031_ = X[401] & Y[401];
assign S[401] = _3030_ ^ _3029_;
assign _3033_ = _3030_ & _3029_;
assign _3034_ = _3031_ | _3033_;
assign _3035_ = X[402] ^ Y[402];
assign _3036_ = X[402] & Y[402];
assign S[402] = _3035_ ^ _3034_;
assign _3038_ = _3035_ & _3034_;
assign _3039_ = _3036_ | _3038_;
assign _3040_ = X[403] ^ Y[403];
assign _3041_ = X[403] & Y[403];
assign S[403] = _3040_ ^ _3039_;
assign _3043_ = _3040_ & _3039_;
assign _3044_ = _3041_ | _3043_;
assign _3045_ = X[404] ^ Y[404];
assign _3046_ = X[404] & Y[404];
assign S[404] = _3045_ ^ _3044_;
assign _3048_ = _3045_ & _3044_;
assign _3049_ = _3046_ | _3048_;
assign _3050_ = X[405] ^ Y[405];
assign _3051_ = X[405] & Y[405];
assign S[405] = _3050_ ^ _3049_;
assign _3053_ = _3050_ & _3049_;
assign _3054_ = _3051_ | _3053_;
assign _3055_ = X[406] ^ Y[406];
assign _3056_ = X[406] & Y[406];
assign S[406] = _3055_ ^ _3054_;
assign _3058_ = _3055_ & _3054_;
assign _3059_ = _3056_ | _3058_;
assign _3060_ = X[407] ^ Y[407];
assign _3061_ = X[407] & Y[407];
assign S[407] = _3060_ ^ _3059_;
assign _3063_ = _3060_ & _3059_;
assign _3064_ = _3061_ | _3063_;
assign _3065_ = X[408] ^ Y[408];
assign _3066_ = X[408] & Y[408];
assign S[408] = _3065_ ^ _3064_;
assign _3068_ = _3065_ & _3064_;
assign _3069_ = _3066_ | _3068_;
assign _3070_ = X[409] ^ Y[409];
assign _3071_ = X[409] & Y[409];
assign S[409] = _3070_ ^ _3069_;
assign _3073_ = _3070_ & _3069_;
assign _3074_ = _3071_ | _3073_;
assign _3075_ = X[410] ^ Y[410];
assign _3076_ = X[410] & Y[410];
assign S[410] = _3075_ ^ _3074_;
assign _3078_ = _3075_ & _3074_;
assign _3079_ = _3076_ | _3078_;
assign _3080_ = X[411] ^ Y[411];
assign _3081_ = X[411] & Y[411];
assign S[411] = _3080_ ^ _3079_;
assign _3083_ = _3080_ & _3079_;
assign _3084_ = _3081_ | _3083_;
assign _3085_ = X[412] ^ Y[412];
assign _3086_ = X[412] & Y[412];
assign S[412] = _3085_ ^ _3084_;
assign _3088_ = _3085_ & _3084_;
assign _3089_ = _3086_ | _3088_;
assign _3090_ = X[413] ^ Y[413];
assign _3091_ = X[413] & Y[413];
assign S[413] = _3090_ ^ _3089_;
assign _3093_ = _3090_ & _3089_;
assign _3094_ = _3091_ | _3093_;
assign _3095_ = X[414] ^ Y[414];
assign _3096_ = X[414] & Y[414];
assign S[414] = _3095_ ^ _3094_;
assign _3098_ = _3095_ & _3094_;
assign _3099_ = _3096_ | _3098_;
assign _3100_ = X[415] ^ Y[415];
assign _3101_ = X[415] & Y[415];
assign S[415] = _3100_ ^ _3099_;
assign _3103_ = _3100_ & _3099_;
assign _3104_ = _3101_ | _3103_;
assign _3105_ = X[416] ^ Y[416];
assign _3106_ = X[416] & Y[416];
assign S[416] = _3105_ ^ _3104_;
assign _3108_ = _3105_ & _3104_;
assign _3109_ = _3106_ | _3108_;
assign _3110_ = X[417] ^ Y[417];
assign _3111_ = X[417] & Y[417];
assign S[417] = _3110_ ^ _3109_;
assign _3113_ = _3110_ & _3109_;
assign _3114_ = _3111_ | _3113_;
assign _3115_ = X[418] ^ Y[418];
assign _3116_ = X[418] & Y[418];
assign S[418] = _3115_ ^ _3114_;
assign _3118_ = _3115_ & _3114_;
assign _3119_ = _3116_ | _3118_;
assign _3120_ = X[419] ^ Y[419];
assign _3121_ = X[419] & Y[419];
assign S[419] = _3120_ ^ _3119_;
assign _3123_ = _3120_ & _3119_;
assign _3124_ = _3121_ | _3123_;
assign _3125_ = X[420] ^ Y[420];
assign _3126_ = X[420] & Y[420];
assign S[420] = _3125_ ^ _3124_;
assign _3128_ = _3125_ & _3124_;
assign _3129_ = _3126_ | _3128_;
assign _3130_ = X[421] ^ Y[421];
assign _3131_ = X[421] & Y[421];
assign S[421] = _3130_ ^ _3129_;
assign _3133_ = _3130_ & _3129_;
assign _3134_ = _3131_ | _3133_;
assign _3135_ = X[422] ^ Y[422];
assign _3136_ = X[422] & Y[422];
assign S[422] = _3135_ ^ _3134_;
assign _3138_ = _3135_ & _3134_;
assign _3139_ = _3136_ | _3138_;
assign _3140_ = X[423] ^ Y[423];
assign _3141_ = X[423] & Y[423];
assign S[423] = _3140_ ^ _3139_;
assign _3143_ = _3140_ & _3139_;
assign _3144_ = _3141_ | _3143_;
assign _3145_ = X[424] ^ Y[424];
assign _3146_ = X[424] & Y[424];
assign S[424] = _3145_ ^ _3144_;
assign _3148_ = _3145_ & _3144_;
assign _3149_ = _3146_ | _3148_;
assign _3150_ = X[425] ^ Y[425];
assign _3151_ = X[425] & Y[425];
assign S[425] = _3150_ ^ _3149_;
assign _3153_ = _3150_ & _3149_;
assign _3154_ = _3151_ | _3153_;
assign _3155_ = X[426] ^ Y[426];
assign _3156_ = X[426] & Y[426];
assign S[426] = _3155_ ^ _3154_;
assign _3158_ = _3155_ & _3154_;
assign _3159_ = _3156_ | _3158_;
assign _3160_ = X[427] ^ Y[427];
assign _3161_ = X[427] & Y[427];
assign S[427] = _3160_ ^ _3159_;
assign _3163_ = _3160_ & _3159_;
assign _3164_ = _3161_ | _3163_;
assign _3165_ = X[428] ^ Y[428];
assign _3166_ = X[428] & Y[428];
assign S[428] = _3165_ ^ _3164_;
assign _3168_ = _3165_ & _3164_;
assign _3169_ = _3166_ | _3168_;
assign _3170_ = X[429] ^ Y[429];
assign _3171_ = X[429] & Y[429];
assign S[429] = _3170_ ^ _3169_;
assign _3173_ = _3170_ & _3169_;
assign _3174_ = _3171_ | _3173_;
assign _3175_ = X[430] ^ Y[430];
assign _3176_ = X[430] & Y[430];
assign S[430] = _3175_ ^ _3174_;
assign _3178_ = _3175_ & _3174_;
assign _3179_ = _3176_ | _3178_;
assign _3180_ = X[431] ^ Y[431];
assign _3181_ = X[431] & Y[431];
assign S[431] = _3180_ ^ _3179_;
assign _3183_ = _3180_ & _3179_;
assign _3184_ = _3181_ | _3183_;
assign _3185_ = X[432] ^ Y[432];
assign _3186_ = X[432] & Y[432];
assign S[432] = _3185_ ^ _3184_;
assign _3188_ = _3185_ & _3184_;
assign _3189_ = _3186_ | _3188_;
assign _3190_ = X[433] ^ Y[433];
assign _3191_ = X[433] & Y[433];
assign S[433] = _3190_ ^ _3189_;
assign _3193_ = _3190_ & _3189_;
assign _3194_ = _3191_ | _3193_;
assign _3195_ = X[434] ^ Y[434];
assign _3196_ = X[434] & Y[434];
assign S[434] = _3195_ ^ _3194_;
assign _3198_ = _3195_ & _3194_;
assign _3199_ = _3196_ | _3198_;
assign _3200_ = X[435] ^ Y[435];
assign _3201_ = X[435] & Y[435];
assign S[435] = _3200_ ^ _3199_;
assign _3203_ = _3200_ & _3199_;
assign _3204_ = _3201_ | _3203_;
assign _3205_ = X[436] ^ Y[436];
assign _3206_ = X[436] & Y[436];
assign S[436] = _3205_ ^ _3204_;
assign _3208_ = _3205_ & _3204_;
assign _3209_ = _3206_ | _3208_;
assign _3210_ = X[437] ^ Y[437];
assign _3211_ = X[437] & Y[437];
assign S[437] = _3210_ ^ _3209_;
assign _3213_ = _3210_ & _3209_;
assign _3214_ = _3211_ | _3213_;
assign _3215_ = X[438] ^ Y[438];
assign _3216_ = X[438] & Y[438];
assign S[438] = _3215_ ^ _3214_;
assign _3218_ = _3215_ & _3214_;
assign _3219_ = _3216_ | _3218_;
assign _3220_ = X[439] ^ Y[439];
assign _3221_ = X[439] & Y[439];
assign S[439] = _3220_ ^ _3219_;
assign _3223_ = _3220_ & _3219_;
assign _3224_ = _3221_ | _3223_;
assign _3225_ = X[440] ^ Y[440];
assign _3226_ = X[440] & Y[440];
assign S[440] = _3225_ ^ _3224_;
assign _3228_ = _3225_ & _3224_;
assign _3229_ = _3226_ | _3228_;
assign _3230_ = X[441] ^ Y[441];
assign _3231_ = X[441] & Y[441];
assign S[441] = _3230_ ^ _3229_;
assign _3233_ = _3230_ & _3229_;
assign _3234_ = _3231_ | _3233_;
assign _3235_ = X[442] ^ Y[442];
assign _3236_ = X[442] & Y[442];
assign S[442] = _3235_ ^ _3234_;
assign _3238_ = _3235_ & _3234_;
assign _3239_ = _3236_ | _3238_;
assign _3240_ = X[443] ^ Y[443];
assign _3241_ = X[443] & Y[443];
assign S[443] = _3240_ ^ _3239_;
assign _3243_ = _3240_ & _3239_;
assign _3244_ = _3241_ | _3243_;
assign _3245_ = X[444] ^ Y[444];
assign _3246_ = X[444] & Y[444];
assign S[444] = _3245_ ^ _3244_;
assign _3248_ = _3245_ & _3244_;
assign _3249_ = _3246_ | _3248_;
assign _3250_ = X[445] ^ Y[445];
assign _3251_ = X[445] & Y[445];
assign S[445] = _3250_ ^ _3249_;
assign _3253_ = _3250_ & _3249_;
assign _3254_ = _3251_ | _3253_;
assign _3255_ = X[446] ^ Y[446];
assign _3256_ = X[446] & Y[446];
assign S[446] = _3255_ ^ _3254_;
assign _3258_ = _3255_ & _3254_;
assign _3259_ = _3256_ | _3258_;
assign _3260_ = X[447] ^ Y[447];
assign _3261_ = X[447] & Y[447];
assign S[447] = _3260_ ^ _3259_;
assign _3263_ = _3260_ & _3259_;
assign _3264_ = _3261_ | _3263_;
assign _3265_ = X[448] ^ Y[448];
assign _3266_ = X[448] & Y[448];
assign S[448] = _3265_ ^ _3264_;
assign _3268_ = _3265_ & _3264_;
assign _3269_ = _3266_ | _3268_;
assign _3270_ = X[449] ^ Y[449];
assign _3271_ = X[449] & Y[449];
assign S[449] = _3270_ ^ _3269_;
assign _3273_ = _3270_ & _3269_;
assign _3274_ = _3271_ | _3273_;
assign _3275_ = X[450] ^ Y[450];
assign _3276_ = X[450] & Y[450];
assign S[450] = _3275_ ^ _3274_;
assign _3278_ = _3275_ & _3274_;
assign _3279_ = _3276_ | _3278_;
assign _3280_ = X[451] ^ Y[451];
assign _3281_ = X[451] & Y[451];
assign S[451] = _3280_ ^ _3279_;
assign _3283_ = _3280_ & _3279_;
assign _3284_ = _3281_ | _3283_;
assign _3285_ = X[452] ^ Y[452];
assign _3286_ = X[452] & Y[452];
assign S[452] = _3285_ ^ _3284_;
assign _3288_ = _3285_ & _3284_;
assign _3289_ = _3286_ | _3288_;
assign _3290_ = X[453] ^ Y[453];
assign _3291_ = X[453] & Y[453];
assign S[453] = _3290_ ^ _3289_;
assign _3293_ = _3290_ & _3289_;
assign _3294_ = _3291_ | _3293_;
assign _3295_ = X[454] ^ Y[454];
assign _3296_ = X[454] & Y[454];
assign S[454] = _3295_ ^ _3294_;
assign _3298_ = _3295_ & _3294_;
assign _3299_ = _3296_ | _3298_;
assign _3300_ = X[455] ^ Y[455];
assign _3301_ = X[455] & Y[455];
assign S[455] = _3300_ ^ _3299_;
assign _3303_ = _3300_ & _3299_;
assign _3304_ = _3301_ | _3303_;
assign _3305_ = X[456] ^ Y[456];
assign _3306_ = X[456] & Y[456];
assign S[456] = _3305_ ^ _3304_;
assign _3308_ = _3305_ & _3304_;
assign _3309_ = _3306_ | _3308_;
assign _3310_ = X[457] ^ Y[457];
assign _3311_ = X[457] & Y[457];
assign S[457] = _3310_ ^ _3309_;
assign _3313_ = _3310_ & _3309_;
assign _3314_ = _3311_ | _3313_;
assign _3315_ = X[458] ^ Y[458];
assign _3316_ = X[458] & Y[458];
assign S[458] = _3315_ ^ _3314_;
assign _3318_ = _3315_ & _3314_;
assign _3319_ = _3316_ | _3318_;
assign _3320_ = X[459] ^ Y[459];
assign _3321_ = X[459] & Y[459];
assign S[459] = _3320_ ^ _3319_;
assign _3323_ = _3320_ & _3319_;
assign _3324_ = _3321_ | _3323_;
assign _3325_ = X[460] ^ Y[460];
assign _3326_ = X[460] & Y[460];
assign S[460] = _3325_ ^ _3324_;
assign _3328_ = _3325_ & _3324_;
assign _3329_ = _3326_ | _3328_;
assign _3330_ = X[461] ^ Y[461];
assign _3331_ = X[461] & Y[461];
assign S[461] = _3330_ ^ _3329_;
assign _3333_ = _3330_ & _3329_;
assign _3334_ = _3331_ | _3333_;
assign _3335_ = X[462] ^ Y[462];
assign _3336_ = X[462] & Y[462];
assign S[462] = _3335_ ^ _3334_;
assign _3338_ = _3335_ & _3334_;
assign _3339_ = _3336_ | _3338_;
assign _3340_ = X[463] ^ Y[463];
assign _3341_ = X[463] & Y[463];
assign S[463] = _3340_ ^ _3339_;
assign _3343_ = _3340_ & _3339_;
assign _3344_ = _3341_ | _3343_;
assign _3345_ = X[464] ^ Y[464];
assign _3346_ = X[464] & Y[464];
assign S[464] = _3345_ ^ _3344_;
assign _3348_ = _3345_ & _3344_;
assign _3349_ = _3346_ | _3348_;
assign _3350_ = X[465] ^ Y[465];
assign _3351_ = X[465] & Y[465];
assign S[465] = _3350_ ^ _3349_;
assign _3353_ = _3350_ & _3349_;
assign _3354_ = _3351_ | _3353_;
assign _3355_ = X[466] ^ Y[466];
assign _3356_ = X[466] & Y[466];
assign S[466] = _3355_ ^ _3354_;
assign _3358_ = _3355_ & _3354_;
assign _3359_ = _3356_ | _3358_;
assign _3360_ = X[467] ^ Y[467];
assign _3361_ = X[467] & Y[467];
assign S[467] = _3360_ ^ _3359_;
assign _3363_ = _3360_ & _3359_;
assign _3364_ = _3361_ | _3363_;
assign _3365_ = X[468] ^ Y[468];
assign _3366_ = X[468] & Y[468];
assign S[468] = _3365_ ^ _3364_;
assign _3368_ = _3365_ & _3364_;
assign _3369_ = _3366_ | _3368_;
assign _3370_ = X[469] ^ Y[469];
assign _3371_ = X[469] & Y[469];
assign S[469] = _3370_ ^ _3369_;
assign _3373_ = _3370_ & _3369_;
assign _3374_ = _3371_ | _3373_;
assign _3375_ = X[470] ^ Y[470];
assign _3376_ = X[470] & Y[470];
assign S[470] = _3375_ ^ _3374_;
assign _3378_ = _3375_ & _3374_;
assign _3379_ = _3376_ | _3378_;
assign _3380_ = X[471] ^ Y[471];
assign _3381_ = X[471] & Y[471];
assign S[471] = _3380_ ^ _3379_;
assign _3383_ = _3380_ & _3379_;
assign _3384_ = _3381_ | _3383_;
assign _3385_ = X[472] ^ Y[472];
assign _3386_ = X[472] & Y[472];
assign S[472] = _3385_ ^ _3384_;
assign _3388_ = _3385_ & _3384_;
assign _3389_ = _3386_ | _3388_;
assign _3390_ = X[473] ^ Y[473];
assign _3391_ = X[473] & Y[473];
assign S[473] = _3390_ ^ _3389_;
assign _3393_ = _3390_ & _3389_;
assign _3394_ = _3391_ | _3393_;
assign _3395_ = X[474] ^ Y[474];
assign _3396_ = X[474] & Y[474];
assign S[474] = _3395_ ^ _3394_;
assign _3398_ = _3395_ & _3394_;
assign _3399_ = _3396_ | _3398_;
assign _3400_ = X[475] ^ Y[475];
assign _3401_ = X[475] & Y[475];
assign S[475] = _3400_ ^ _3399_;
assign _3403_ = _3400_ & _3399_;
assign _3404_ = _3401_ | _3403_;
assign _3405_ = X[476] ^ Y[476];
assign _3406_ = X[476] & Y[476];
assign S[476] = _3405_ ^ _3404_;
assign _3408_ = _3405_ & _3404_;
assign _3409_ = _3406_ | _3408_;
assign _3410_ = X[477] ^ Y[477];
assign _3411_ = X[477] & Y[477];
assign S[477] = _3410_ ^ _3409_;
assign _3413_ = _3410_ & _3409_;
assign _3414_ = _3411_ | _3413_;
assign _3415_ = X[478] ^ Y[478];
assign _3416_ = X[478] & Y[478];
assign S[478] = _3415_ ^ _3414_;
assign _3418_ = _3415_ & _3414_;
assign _3419_ = _3416_ | _3418_;
assign _3420_ = X[479] ^ Y[479];
assign _3421_ = X[479] & Y[479];
assign S[479] = _3420_ ^ _3419_;
assign _3423_ = _3420_ & _3419_;
assign _3424_ = _3421_ | _3423_;
assign _3425_ = X[480] ^ Y[480];
assign _3426_ = X[480] & Y[480];
assign S[480] = _3425_ ^ _3424_;
assign _3428_ = _3425_ & _3424_;
assign _3429_ = _3426_ | _3428_;
assign _3430_ = X[481] ^ Y[481];
assign _3431_ = X[481] & Y[481];
assign S[481] = _3430_ ^ _3429_;
assign _3433_ = _3430_ & _3429_;
assign _3434_ = _3431_ | _3433_;
assign _3435_ = X[482] ^ Y[482];
assign _3436_ = X[482] & Y[482];
assign S[482] = _3435_ ^ _3434_;
assign _3438_ = _3435_ & _3434_;
assign _3439_ = _3436_ | _3438_;
assign _3440_ = X[483] ^ Y[483];
assign _3441_ = X[483] & Y[483];
assign S[483] = _3440_ ^ _3439_;
assign _3443_ = _3440_ & _3439_;
assign _3444_ = _3441_ | _3443_;
assign _3445_ = X[484] ^ Y[484];
assign _3446_ = X[484] & Y[484];
assign S[484] = _3445_ ^ _3444_;
assign _3448_ = _3445_ & _3444_;
assign _3449_ = _3446_ | _3448_;
assign _3450_ = X[485] ^ Y[485];
assign _3451_ = X[485] & Y[485];
assign S[485] = _3450_ ^ _3449_;
assign _3453_ = _3450_ & _3449_;
assign _3454_ = _3451_ | _3453_;
assign _3455_ = X[486] ^ Y[486];
assign _3456_ = X[486] & Y[486];
assign S[486] = _3455_ ^ _3454_;
assign _3458_ = _3455_ & _3454_;
assign _3459_ = _3456_ | _3458_;
assign _3460_ = X[487] ^ Y[487];
assign _3461_ = X[487] & Y[487];
assign S[487] = _3460_ ^ _3459_;
assign _3463_ = _3460_ & _3459_;
assign _3464_ = _3461_ | _3463_;
assign _3465_ = X[488] ^ Y[488];
assign _3466_ = X[488] & Y[488];
assign S[488] = _3465_ ^ _3464_;
assign _3468_ = _3465_ & _3464_;
assign _3469_ = _3466_ | _3468_;
assign _3470_ = X[489] ^ Y[489];
assign _3471_ = X[489] & Y[489];
assign S[489] = _3470_ ^ _3469_;
assign _3473_ = _3470_ & _3469_;
assign _3474_ = _3471_ | _3473_;
assign _3475_ = X[490] ^ Y[490];
assign _3476_ = X[490] & Y[490];
assign S[490] = _3475_ ^ _3474_;
assign _3478_ = _3475_ & _3474_;
assign _3479_ = _3476_ | _3478_;
assign _3480_ = X[491] ^ Y[491];
assign _3481_ = X[491] & Y[491];
assign S[491] = _3480_ ^ _3479_;
assign _3483_ = _3480_ & _3479_;
assign _3484_ = _3481_ | _3483_;
assign _3485_ = X[492] ^ Y[492];
assign _3486_ = X[492] & Y[492];
assign S[492] = _3485_ ^ _3484_;
assign _3488_ = _3485_ & _3484_;
assign _3489_ = _3486_ | _3488_;
assign _3490_ = X[493] ^ Y[493];
assign _3491_ = X[493] & Y[493];
assign S[493] = _3490_ ^ _3489_;
assign _3493_ = _3490_ & _3489_;
assign _3494_ = _3491_ | _3493_;
assign _3495_ = X[494] ^ Y[494];
assign _3496_ = X[494] & Y[494];
assign S[494] = _3495_ ^ _3494_;
assign _3498_ = _3495_ & _3494_;
assign _3499_ = _3496_ | _3498_;
assign _3500_ = X[495] ^ Y[495];
assign _3501_ = X[495] & Y[495];
assign S[495] = _3500_ ^ _3499_;
assign _3503_ = _3500_ & _3499_;
assign _3504_ = _3501_ | _3503_;
assign _3505_ = X[496] ^ Y[496];
assign _3506_ = X[496] & Y[496];
assign S[496] = _3505_ ^ _3504_;
assign _3508_ = _3505_ & _3504_;
assign _3509_ = _3506_ | _3508_;
assign _3510_ = X[497] ^ Y[497];
assign _3511_ = X[497] & Y[497];
assign S[497] = _3510_ ^ _3509_;
assign _3513_ = _3510_ & _3509_;
assign _3514_ = _3511_ | _3513_;
assign _3515_ = X[498] ^ Y[498];
assign _3516_ = X[498] & Y[498];
assign S[498] = _3515_ ^ _3514_;
assign _3518_ = _3515_ & _3514_;
assign _3519_ = _3516_ | _3518_;
assign _3520_ = X[499] ^ Y[499];
assign _3521_ = X[499] & Y[499];
assign S[499] = _3520_ ^ _3519_;
assign _3523_ = _3520_ & _3519_;
assign _3524_ = _3521_ | _3523_;
assign _3525_ = X[500] ^ Y[500];
assign _3526_ = X[500] & Y[500];
assign S[500] = _3525_ ^ _3524_;
assign _3528_ = _3525_ & _3524_;
assign _3529_ = _3526_ | _3528_;
assign _3530_ = X[501] ^ Y[501];
assign _3531_ = X[501] & Y[501];
assign S[501] = _3530_ ^ _3529_;
assign _3533_ = _3530_ & _3529_;
assign _3534_ = _3531_ | _3533_;
assign _3535_ = X[502] ^ Y[502];
assign _3536_ = X[502] & Y[502];
assign S[502] = _3535_ ^ _3534_;
assign _3538_ = _3535_ & _3534_;
assign _3539_ = _3536_ | _3538_;
assign _3540_ = X[503] ^ Y[503];
assign _3541_ = X[503] & Y[503];
assign S[503] = _3540_ ^ _3539_;
assign _3543_ = _3540_ & _3539_;
assign _3544_ = _3541_ | _3543_;
assign _3545_ = X[504] ^ Y[504];
assign _3546_ = X[504] & Y[504];
assign S[504] = _3545_ ^ _3544_;
assign _3548_ = _3545_ & _3544_;
assign _3549_ = _3546_ | _3548_;
assign _3550_ = X[505] ^ Y[505];
assign _3551_ = X[505] & Y[505];
assign S[505] = _3550_ ^ _3549_;
assign _3553_ = _3550_ & _3549_;
assign _3554_ = _3551_ | _3553_;
assign _3555_ = X[506] ^ Y[506];
assign _3556_ = X[506] & Y[506];
assign S[506] = _3555_ ^ _3554_;
assign _3558_ = _3555_ & _3554_;
assign _3559_ = _3556_ | _3558_;
assign _3560_ = X[507] ^ Y[507];
assign _3561_ = X[507] & Y[507];
assign S[507] = _3560_ ^ _3559_;
assign _3563_ = _3560_ & _3559_;
assign _3564_ = _3561_ | _3563_;
assign _3565_ = X[508] ^ Y[508];
assign _3566_ = X[508] & Y[508];
assign S[508] = _3565_ ^ _3564_;
assign _3568_ = _3565_ & _3564_;
assign _3569_ = _3566_ | _3568_;
assign _3570_ = X[509] ^ Y[509];
assign _3571_ = X[509] & Y[509];
assign S[509] = _3570_ ^ _3569_;
assign _3573_ = _3570_ & _3569_;
assign _3574_ = _3571_ | _3573_;
assign _3575_ = X[510] ^ Y[510];
assign _3576_ = X[510] & Y[510];
assign S[510] = _3575_ ^ _3574_;
assign _3578_ = _3575_ & _3574_;
assign _3579_ = _3576_ | _3578_;
assign _3580_ = X[511] ^ Y[511];
assign _3581_ = X[511] & Y[511];
assign S[511] = _3580_ ^ _3579_;
assign _3583_ = _3580_ & _3579_;
assign S[512] = _3581_ | _3583_;
endmodule